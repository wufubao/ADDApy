assign q[0]= 16'h389;
assign q[1]= 16'h669;
assign q[2]= 16'h901;
assign q[3]= 16'hb32;
assign q[4]= 16'hcde;
assign q[5]= 16'hdec;
assign q[6]= 16'he49;
assign q[7]= 16'hde7;
assign q[8]= 16'hcc2;
assign q[9]= 16'hada;
assign q[10]= 16'h83a;
assign q[11]= 16'h4f0;
assign q[12]= 16'h115;
assign q[13]= 16'hfcc7;
assign q[14]= 16'hf826;
assign q[15]= 16'hf359;
assign q[16]= 16'hee89;
assign q[17]= 16'he9e1;
assign q[18]= 16'he58a;
assign q[19]= 16'he1ab;
assign q[20]= 16'hde69;
assign q[21]= 16'hdbe4;
assign q[22]= 16'hda36;
assign q[23]= 16'hd973;
assign q[24]= 16'hd9a7;
assign q[25]= 16'hdad6;
assign q[26]= 16'hdcfd;
assign q[27]= 16'he012;
assign q[28]= 16'he401;
assign q[29]= 16'he8b1;
assign q[30]= 16'hee04;
assign q[31]= 16'hf3d5;
assign q[32]= 16'hf9fe;
assign q[33]= 16'h52;
assign q[34]= 16'h6aa;
assign q[35]= 16'hcda;
assign q[36]= 16'h12b8;
assign q[37]= 16'h1820;
assign q[38]= 16'h1cef;
assign q[39]= 16'h2107;
assign q[40]= 16'h2451;
assign q[41]= 16'h26bb;
assign q[42]= 16'h2839;
assign q[43]= 16'h28c7;
assign q[44]= 16'h2865;
assign q[45]= 16'h271b;
assign q[46]= 16'h24f6;
assign q[47]= 16'h2206;
assign q[48]= 16'h1e62;
assign q[49]= 16'h1a22;
assign q[50]= 16'h1561;
assign q[51]= 16'h103d;
assign q[52]= 16'had3;
assign q[53]= 16'h540;
assign q[54]= 16'hffa1;
assign q[55]= 16'hfa10;
assign q[56]= 16'hf4a6;
assign q[57]= 16'hef7a;
assign q[58]= 16'hea9e;
assign q[59]= 16'he624;
assign q[60]= 16'he218;
assign q[61]= 16'hde84;
assign q[62]= 16'hdb70;
assign q[63]= 16'hd8df;
assign q[64]= 16'hd6d1;
assign q[65]= 16'hd547;
assign q[66]= 16'hd43d;
assign q[67]= 16'hd3ac;
assign q[68]= 16'hd38e;
assign q[69]= 16'hd3da;
assign q[70]= 16'hd487;
assign q[71]= 16'hd589;
assign q[72]= 16'hd6d7;
assign q[73]= 16'hd862;
assign q[74]= 16'hda20;
assign q[75]= 16'hdc04;
assign q[76]= 16'hde01;
assign q[77]= 16'he00a;
assign q[78]= 16'he213;
assign q[79]= 16'he40f;
assign q[80]= 16'he5f3;
assign q[81]= 16'he7b4;
assign q[82]= 16'he948;
assign q[83]= 16'heaa4;
assign q[84]= 16'hebc1;
assign q[85]= 16'hec98;
assign q[86]= 16'hed24;
assign q[87]= 16'hed61;
assign q[88]= 16'hed4d;
assign q[89]= 16'hecea;
assign q[90]= 16'hec38;
assign q[91]= 16'heb3e;
assign q[92]= 16'hea01;
assign q[93]= 16'he88b;
assign q[94]= 16'he6e5;
assign q[95]= 16'he51d;
assign q[96]= 16'he33f;
assign q[97]= 16'he15c;
assign q[98]= 16'hdf82;
assign q[99]= 16'hddc2;
assign q[100]= 16'hdc2c;
assign q[101]= 16'hdacf;
assign q[102]= 16'hd9bb;
assign q[103]= 16'hd8fd;
assign q[104]= 16'hd8a1;
assign q[105]= 16'hd8b2;
assign q[106]= 16'hd938;
assign q[107]= 16'hda38;
assign q[108]= 16'hdbb6;
assign q[109]= 16'hddb3;
assign q[110]= 16'he02b;
assign q[111]= 16'he31b;
assign q[112]= 16'he67b;
assign q[113]= 16'hea41;
assign q[114]= 16'hee63;
assign q[115]= 16'hf2d1;
assign q[116]= 16'hf77d;
assign q[117]= 16'hfc56;
assign q[118]= 16'h14a;
assign q[119]= 16'h649;
assign q[120]= 16'hb3e;
assign q[121]= 16'h1019;
assign q[122]= 16'h14c7;
assign q[123]= 16'h1936;
assign q[124]= 16'h1d56;
assign q[125]= 16'h2118;
assign q[126]= 16'h246e;
assign q[127]= 16'h274a;
assign q[128]= 16'h29a3;
assign q[129]= 16'h2b6f;
assign q[130]= 16'h2ca7;
assign q[131]= 16'h2d46;
assign q[132]= 16'h2d49;
assign q[133]= 16'h2cae;
assign q[134]= 16'h2b77;
assign q[135]= 16'h29a6;
assign q[136]= 16'h2740;
assign q[137]= 16'h244e;
assign q[138]= 16'h20d7;
assign q[139]= 16'h1ce6;
assign q[140]= 16'h1889;
assign q[141]= 16'h13cd;
assign q[142]= 16'hec1;
assign q[143]= 16'h977;
assign q[144]= 16'h400;
assign q[145]= 16'hfe6e;
assign q[146]= 16'hf8d3;
assign q[147]= 16'hf343;
assign q[148]= 16'hedcf;
assign q[149]= 16'he889;
assign q[150]= 16'he383;
assign q[151]= 16'hdecc;
assign q[152]= 16'hda72;
assign q[153]= 16'hd683;
assign q[154]= 16'hd307;
assign q[155]= 16'hd009;
assign q[156]= 16'hcd8d;
assign q[157]= 16'hcb99;
assign q[158]= 16'hca2d;
assign q[159]= 16'hc949;
assign q[160]= 16'hc8eb;
assign q[161]= 16'hc90c;
assign q[162]= 16'hc9a8;
assign q[163]= 16'hcab6;
assign q[164]= 16'hcc2c;
assign q[165]= 16'hce02;
assign q[166]= 16'hd02c;
assign q[167]= 16'hd29f;
assign q[168]= 16'hd551;
assign q[169]= 16'hd839;
assign q[170]= 16'hdb4b;
assign q[171]= 16'hde7f;
assign q[172]= 16'he1cd;
assign q[173]= 16'he52e;
assign q[174]= 16'he89c;
assign q[175]= 16'hec12;
assign q[176]= 16'hef8d;
assign q[177]= 16'hf30a;
assign q[178]= 16'hf685;
assign q[179]= 16'hf9fe;
assign q[180]= 16'hfd73;
assign q[181]= 16'he1;
assign q[182]= 16'h449;
assign q[183]= 16'h7a7;
assign q[184]= 16'hafa;
assign q[185]= 16'he3e;
assign q[186]= 16'h1170;
assign q[187]= 16'h148b;
assign q[188]= 16'h178a;
assign q[189]= 16'h1a68;
assign q[190]= 16'h1d1d;
assign q[191]= 16'h1fa3;
assign q[192]= 16'h21f4;
assign q[193]= 16'h2408;
assign q[194]= 16'h25da;
assign q[195]= 16'h2762;
assign q[196]= 16'h289d;
assign q[197]= 16'h2985;
assign q[198]= 16'h2a19;
assign q[199]= 16'h2a57;
assign q[200]= 16'h2a40;
assign q[201]= 16'h29d5;
assign q[202]= 16'h291b;
assign q[203]= 16'h2815;
assign q[204]= 16'h26cc;
assign q[205]= 16'h2547;
assign q[206]= 16'h2390;
assign q[207]= 16'h21b0;
assign q[208]= 16'h1fb3;
assign q[209]= 16'h1da4;
assign q[210]= 16'h1b8d;
assign q[211]= 16'h197a;
assign q[212]= 16'h1775;
assign q[213]= 16'h1587;
assign q[214]= 16'h13b8;
assign q[215]= 16'h1210;
assign q[216]= 16'h1095;
assign q[217]= 16'hf4a;
assign q[218]= 16'he32;
assign q[219]= 16'hd4e;
assign q[220]= 16'hc9f;
assign q[221]= 16'hc21;
assign q[222]= 16'hbd3;
assign q[223]= 16'hbb1;
assign q[224]= 16'hbb6;
assign q[225]= 16'hbdd;
assign q[226]= 16'hc21;
assign q[227]= 16'hc7b;
assign q[228]= 16'hce6;
assign q[229]= 16'hd5d;
assign q[230]= 16'hdda;
assign q[231]= 16'he59;
assign q[232]= 16'hed6;
assign q[233]= 16'hf4c;
assign q[234]= 16'hfb9;
assign q[235]= 16'h1019;
assign q[236]= 16'h106b;
assign q[237]= 16'h10ad;
assign q[238]= 16'h10dc;
assign q[239]= 16'h10f9;
assign q[240]= 16'h1100;
assign q[241]= 16'h10f2;
assign q[242]= 16'h10cd;
assign q[243]= 16'h1090;
assign q[244]= 16'h1039;
assign q[245]= 16'hfc7;
assign q[246]= 16'hf38;
assign q[247]= 16'he8c;
assign q[248]= 16'hdc0;
assign q[249]= 16'hcd5;
assign q[250]= 16'hbc8;
assign q[251]= 16'ha99;
assign q[252]= 16'h948;
assign q[253]= 16'h7d6;
assign q[254]= 16'h644;
assign q[255]= 16'h492;
assign q[256]= 16'h2c4;
assign q[257]= 16'hdc;
assign q[258]= 16'hfedd;
assign q[259]= 16'hfccb;
assign q[260]= 16'hfaab;
assign q[261]= 16'hf87f;
assign q[262]= 16'hf64e;
assign q[263]= 16'hf41c;
assign q[264]= 16'hf1ed;
assign q[265]= 16'hefc4;
assign q[266]= 16'heda6;
assign q[267]= 16'heb96;
assign q[268]= 16'he994;
assign q[269]= 16'he7a5;
assign q[270]= 16'he5c7;
assign q[271]= 16'he3fb;
assign q[272]= 16'he242;
assign q[273]= 16'he099;
assign q[274]= 16'hdf00;
assign q[275]= 16'hdd76;
assign q[276]= 16'hdbf8;
assign q[277]= 16'hda87;
assign q[278]= 16'hd920;
assign q[279]= 16'hd7c3;
assign q[280]= 16'hd672;
assign q[281]= 16'hd52e;
assign q[282]= 16'hd3f7;
assign q[283]= 16'hd2d3;
assign q[284]= 16'hd1c5;
assign q[285]= 16'hd0d1;
assign q[286]= 16'hcffe;
assign q[287]= 16'hcf51;
assign q[288]= 16'hced1;
assign q[289]= 16'hce84;
assign q[290]= 16'hce71;
assign q[291]= 16'hce9c;
assign q[292]= 16'hcf09;
assign q[293]= 16'hcfbd;
assign q[294]= 16'hd0b7;
assign q[295]= 16'hd1f8;
assign q[296]= 16'hd37e;
assign q[297]= 16'hd542;
assign q[298]= 16'hd740;
assign q[299]= 16'hd96e;
assign q[300]= 16'hdbc0;
assign q[301]= 16'hde2c;
assign q[302]= 16'he0a2;
assign q[303]= 16'he314;
assign q[304]= 16'he572;
assign q[305]= 16'he7ac;
assign q[306]= 16'he9b4;
assign q[307]= 16'heb7c;
assign q[308]= 16'hecf6;
assign q[309]= 16'hee18;
assign q[310]= 16'heed9;
assign q[311]= 16'hef35;
assign q[312]= 16'hef28;
assign q[313]= 16'heeb2;
assign q[314]= 16'hedd8;
assign q[315]= 16'heca1;
assign q[316]= 16'heb17;
assign q[317]= 16'he946;
assign q[318]= 16'he73e;
assign q[319]= 16'he50f;
assign q[320]= 16'he2cc;
assign q[321]= 16'he087;
assign q[322]= 16'hde54;
assign q[323]= 16'hdc45;
assign q[324]= 16'hda6a;
assign q[325]= 16'hd8d5;
assign q[326]= 16'hd791;
assign q[327]= 16'hd6a9;
assign q[328]= 16'hd624;
assign q[329]= 16'hd608;
assign q[330]= 16'hd653;
assign q[331]= 16'hd705;
assign q[332]= 16'hd816;
assign q[333]= 16'hd97f;
assign q[334]= 16'hdb33;
assign q[335]= 16'hdd25;
assign q[336]= 16'hdf46;
assign q[337]= 16'he187;
assign q[338]= 16'he3d6;
assign q[339]= 16'he622;
assign q[340]= 16'he85e;
assign q[341]= 16'hea79;
assign q[342]= 16'hec69;
assign q[343]= 16'hee22;
assign q[344]= 16'hef9d;
assign q[345]= 16'hf0d5;
assign q[346]= 16'hf1c8;
assign q[347]= 16'hf278;
assign q[348]= 16'hf2e6;
assign q[349]= 16'hf31a;
assign q[350]= 16'hf31b;
assign q[351]= 16'hf2f4;
assign q[352]= 16'hf2b0;
assign q[353]= 16'hf25b;
assign q[354]= 16'hf201;
assign q[355]= 16'hf1b0;
assign q[356]= 16'hf173;
assign q[357]= 16'hf154;
assign q[358]= 16'hf15e;
assign q[359]= 16'hf198;
assign q[360]= 16'hf207;
assign q[361]= 16'hf2b1;
assign q[362]= 16'hf396;
assign q[363]= 16'hf4b5;
assign q[364]= 16'hf60c;
assign q[365]= 16'hf798;
assign q[366]= 16'hf950;
assign q[367]= 16'hfb2f;
assign q[368]= 16'hfd2b;
assign q[369]= 16'hff3b;
assign q[370]= 16'h154;
assign q[371]= 16'h36f;
assign q[372]= 16'h581;
assign q[373]= 16'h781;
assign q[374]= 16'h966;
assign q[375]= 16'hb2a;
assign q[376]= 16'hcc7;
assign q[377]= 16'he36;
assign q[378]= 16'hf75;
assign q[379]= 16'h1081;
assign q[380]= 16'h115a;
assign q[381]= 16'h11fe;
assign q[382]= 16'h126f;
assign q[383]= 16'h12b0;
assign q[384]= 16'h12c3;
assign q[385]= 16'h12ac;
assign q[386]= 16'h126f;
assign q[387]= 16'h1211;
assign q[388]= 16'h1197;
assign q[389]= 16'h1106;
assign q[390]= 16'h1064;
assign q[391]= 16'hfb7;
assign q[392]= 16'hf03;
assign q[393]= 16'he4f;
assign q[394]= 16'hda0;
assign q[395]= 16'hcfb;
assign q[396]= 16'hc66;
assign q[397]= 16'hbe6;
assign q[398]= 16'hb7e;
assign q[399]= 16'hb35;
assign q[400]= 16'hb0d;
assign q[401]= 16'hb0a;
assign q[402]= 16'hb2f;
assign q[403]= 16'hb7f;
assign q[404]= 16'hbfb;
assign q[405]= 16'hca4;
assign q[406]= 16'hd7a;
assign q[407]= 16'he7d;
assign q[408]= 16'hfac;
assign q[409]= 16'h1102;
assign q[410]= 16'h127e;
assign q[411]= 16'h141a;
assign q[412]= 16'h15d2;
assign q[413]= 16'h17a0;
assign q[414]= 16'h197e;
assign q[415]= 16'h1b66;
assign q[416]= 16'h1d50;
assign q[417]= 16'h1f36;
assign q[418]= 16'h2112;
assign q[419]= 16'h22dc;
assign q[420]= 16'h248f;
assign q[421]= 16'h2627;
assign q[422]= 16'h279e;
assign q[423]= 16'h28f1;
assign q[424]= 16'h2a1e;
assign q[425]= 16'h2b23;
assign q[426]= 16'h2c00;
assign q[427]= 16'h2cb6;
assign q[428]= 16'h2d45;
assign q[429]= 16'h2db0;
assign q[430]= 16'h2df9;
assign q[431]= 16'h2e25;
assign q[432]= 16'h2e36;
assign q[433]= 16'h2e31;
assign q[434]= 16'h2e1b;
assign q[435]= 16'h2df6;
assign q[436]= 16'h2dc7;
assign q[437]= 16'h2d92;
assign q[438]= 16'h2d59;
assign q[439]= 16'h2d20;
assign q[440]= 16'h2ce8;
assign q[441]= 16'h2cb3;
assign q[442]= 16'h2c82;
assign q[443]= 16'h2c56;
assign q[444]= 16'h2c30;
assign q[445]= 16'h2c0e;
assign q[446]= 16'h2bf1;
assign q[447]= 16'h2bd7;
assign q[448]= 16'h2bbf;
assign q[449]= 16'h2ba8;
assign q[450]= 16'h2b90;
assign q[451]= 16'h2b76;
assign q[452]= 16'h2b57;
assign q[453]= 16'h2b30;
assign q[454]= 16'h2b00;
assign q[455]= 16'h2ac2;
assign q[456]= 16'h2a75;
assign q[457]= 16'h2a13;
assign q[458]= 16'h2999;
assign q[459]= 16'h2903;
assign q[460]= 16'h284d;
assign q[461]= 16'h2771;
assign q[462]= 16'h266c;
assign q[463]= 16'h2538;
assign q[464]= 16'h23d2;
assign q[465]= 16'h2236;
assign q[466]= 16'h2062;
assign q[467]= 16'h1e54;
assign q[468]= 16'h1c0c;
assign q[469]= 16'h198a;
assign q[470]= 16'h16d3;
assign q[471]= 16'h13eb;
assign q[472]= 16'h10d9;
assign q[473]= 16'hda5;
assign q[474]= 16'ha5b;
assign q[475]= 16'h708;
assign q[476]= 16'h3ba;
assign q[477]= 16'h81;
assign q[478]= 16'hfd6f;
assign q[479]= 16'hfa93;
assign q[480]= 16'hf800;
assign q[481]= 16'hf5c8;
assign q[482]= 16'hf3fa;
assign q[483]= 16'hf2a4;
assign q[484]= 16'hf1d3;
assign q[485]= 16'hf190;
assign q[486]= 16'hf1e2;
assign q[487]= 16'hf2cb;
assign q[488]= 16'hf44a;
assign q[489]= 16'hf659;
assign q[490]= 16'hf8f0;
assign q[491]= 16'hfc01;
assign q[492]= 16'hff7b;
assign q[493]= 16'h349;
assign q[494]= 16'h755;
assign q[495]= 16'hb85;
assign q[496]= 16'hfbd;
assign q[497]= 16'h13e3;
assign q[498]= 16'h17d9;
assign q[499]= 16'h1b86;
assign q[500]= 16'h1ed0;
assign q[501]= 16'h21a0;
assign q[502]= 16'h23e2;
assign q[503]= 16'h2587;
assign q[504]= 16'h2683;
assign q[505]= 16'h26ce;
assign q[506]= 16'h2666;
assign q[507]= 16'h254d;
assign q[508]= 16'h238b;
assign q[509]= 16'h212a;
assign q[510]= 16'h1e3a;
assign q[511]= 16'h1ace;
assign q[512]= 16'h16fb;
assign q[513]= 16'h12d8;
assign q[514]= 16'he7f;
assign q[515]= 16'ha09;
assign q[516]= 16'h590;
assign q[517]= 16'h12b;
assign q[518]= 16'hfcf3;
assign q[519]= 16'hf8fa;
assign q[520]= 16'hf553;
assign q[521]= 16'hf20d;
assign q[522]= 16'hef34;
assign q[523]= 16'hecd0;
assign q[524]= 16'heae6;
assign q[525]= 16'he977;
assign q[526]= 16'he882;
assign q[527]= 16'he803;
assign q[528]= 16'he7f3;
assign q[529]= 16'he849;
assign q[530]= 16'he8fc;
assign q[531]= 16'hea00;
assign q[532]= 16'heb49;
assign q[533]= 16'heccd;
assign q[534]= 16'hee7f;
assign q[535]= 16'hf054;
assign q[536]= 16'hf242;
assign q[537]= 16'hf43f;
assign q[538]= 16'hf644;
assign q[539]= 16'hf84a;
assign q[540]= 16'hfa4a;
assign q[541]= 16'hfc40;
assign q[542]= 16'hfe28;
assign q[543]= 16'hffff;
assign q[544]= 16'h1c3;
assign q[545]= 16'h372;
assign q[546]= 16'h50b;
assign q[547]= 16'h68d;
assign q[548]= 16'h7f6;
assign q[549]= 16'h947;
assign q[550]= 16'ha7e;
assign q[551]= 16'hb9a;
assign q[552]= 16'hc9a;
assign q[553]= 16'hd7f;
assign q[554]= 16'he46;
assign q[555]= 16'heef;
assign q[556]= 16'hf7b;
assign q[557]= 16'hfe8;
assign q[558]= 16'h1036;
assign q[559]= 16'h1067;
assign q[560]= 16'h107c;
assign q[561]= 16'h1074;
assign q[562]= 16'h1051;
assign q[563]= 16'h1015;
assign q[564]= 16'hfc1;
assign q[565]= 16'hf57;
assign q[566]= 16'hed7;
assign q[567]= 16'he43;
assign q[568]= 16'hd9a;
assign q[569]= 16'hcdd;
assign q[570]= 16'hc0a;
assign q[571]= 16'hb21;
assign q[572]= 16'ha1f;
assign q[573]= 16'h901;
assign q[574]= 16'h7c5;
assign q[575]= 16'h668;
assign q[576]= 16'h4e5;
assign q[577]= 16'h33a;
assign q[578]= 16'h163;
assign q[579]= 16'hff61;
assign q[580]= 16'hfd2f;
assign q[581]= 16'hfad0;
assign q[582]= 16'hf844;
assign q[583]= 16'hf58f;
assign q[584]= 16'hf2b6;
assign q[585]= 16'hefc2;
assign q[586]= 16'hecba;
assign q[587]= 16'he9a9;
assign q[588]= 16'he69d;
assign q[589]= 16'he3a3;
assign q[590]= 16'he0cb;
assign q[591]= 16'hde24;
assign q[592]= 16'hdbbf;
assign q[593]= 16'hd9ac;
assign q[594]= 16'hd7fc;
assign q[595]= 16'hd6bb;
assign q[596]= 16'hd5f9;
assign q[597]= 16'hd5bf;
assign q[598]= 16'hd618;
assign q[599]= 16'hd708;
assign q[600]= 16'hd893;
assign q[601]= 16'hdabb;
assign q[602]= 16'hdd7b;
assign q[603]= 16'he0ce;
assign q[604]= 16'he4ab;
assign q[605]= 16'he906;
assign q[606]= 16'hedd2;
assign q[607]= 16'hf2fd;
assign q[608]= 16'hf877;
assign q[609]= 16'hfe2a;
assign q[610]= 16'h402;
assign q[611]= 16'h9eb;
assign q[612]= 16'hfcf;
assign q[613]= 16'h1599;
assign q[614]= 16'h1b35;
assign q[615]= 16'h2090;
assign q[616]= 16'h2596;
assign q[617]= 16'h2a39;
assign q[618]= 16'h2e68;
assign q[619]= 16'h3216;
assign q[620]= 16'h3539;
assign q[621]= 16'h37c6;
assign q[622]= 16'h39b6;
assign q[623]= 16'h3b04;
assign q[624]= 16'h3bab;
assign q[625]= 16'h3bab;
assign q[626]= 16'h3b02;
assign q[627]= 16'h39b3;
assign q[628]= 16'h37c2;
assign q[629]= 16'h3535;
assign q[630]= 16'h3212;
assign q[631]= 16'h2e63;
assign q[632]= 16'h2a34;
assign q[633]= 16'h2590;
assign q[634]= 16'h2088;
assign q[635]= 16'h1b2a;
assign q[636]= 16'h1589;
assign q[637]= 16'hfb8;
assign q[638]= 16'h9cb;
assign q[639]= 16'h3d7;
assign q[640]= 16'hfdf3;
assign q[641]= 16'hf833;
assign q[642]= 16'hf2ac;
assign q[643]= 16'hed74;
assign q[644]= 16'he89f;
assign q[645]= 16'he43d;
assign q[646]= 16'he05e;
assign q[647]= 16'hdd10;
assign q[648]= 16'hda5d;
assign q[649]= 16'hd84a;
assign q[650]= 16'hd6dc;
assign q[651]= 16'hd612;
assign q[652]= 16'hd5e8;
assign q[653]= 16'hd657;
assign q[654]= 16'hd753;
assign q[655]= 16'hd8cf;
assign q[656]= 16'hdaba;
assign q[657]= 16'hdd02;
assign q[658]= 16'hdf94;
assign q[659]= 16'he25b;
assign q[660]= 16'he543;
assign q[661]= 16'he838;
assign q[662]= 16'heb29;
assign q[663]= 16'hee04;
assign q[664]= 16'hf0bd;
assign q[665]= 16'hf34a;
assign q[666]= 16'hf5a2;
assign q[667]= 16'hf7c3;
assign q[668]= 16'hf9ac;
assign q[669]= 16'hfb60;
assign q[670]= 16'hfce7;
assign q[671]= 16'hfe49;
assign q[672]= 16'hff91;
assign q[673]= 16'hcc;
assign q[674]= 16'h209;
assign q[675]= 16'h355;
assign q[676]= 16'h4bd;
assign q[677]= 16'h64c;
assign q[678]= 16'h80c;
assign q[679]= 16'ha03;
assign q[680]= 16'hc35;
assign q[681]= 16'hea2;
assign q[682]= 16'h1144;
assign q[683]= 16'h1415;
assign q[684]= 16'h1709;
assign q[685]= 16'h1a10;
assign q[686]= 16'h1d18;
assign q[687]= 16'h200e;
assign q[688]= 16'h22db;
assign q[689]= 16'h2569;
assign q[690]= 16'h27a2;
assign q[691]= 16'h2970;
assign q[692]= 16'h2ac1;
assign q[693]= 16'h2b85;
assign q[694]= 16'h2bae;
assign q[695]= 16'h2b34;
assign q[696]= 16'h2a15;
assign q[697]= 16'h2851;
assign q[698]= 16'h25f0;
assign q[699]= 16'h22fe;
assign q[700]= 16'h1f8b;
assign q[701]= 16'h1bae;
assign q[702]= 16'h1780;
assign q[703]= 16'h131e;
assign q[704]= 16'hea6;
assign q[705]= 16'ha39;
assign q[706]= 16'h5f6;
assign q[707]= 16'h1fe;
assign q[708]= 16'hfe6f;
assign q[709]= 16'hfb62;
assign q[710]= 16'hf8ee;
assign q[711]= 16'hf727;
assign q[712]= 16'hf61a;
assign q[713]= 16'hf5cf;
assign q[714]= 16'hf649;
assign q[715]= 16'hf784;
assign q[716]= 16'hf977;
assign q[717]= 16'hfc15;
assign q[718]= 16'hff4a;
assign q[719]= 16'h300;
assign q[720]= 16'h71e;
assign q[721]= 16'hb87;
assign q[722]= 16'h101d;
assign q[723]= 16'h14c4;
assign q[724]= 16'h195e;
assign q[725]= 16'h1dcf;
assign q[726]= 16'h21ff;
assign q[727]= 16'h25d7;
assign q[728]= 16'h2946;
assign q[729]= 16'h2c3d;
assign q[730]= 16'h2eb3;
assign q[731]= 16'h30a4;
assign q[732]= 16'h320f;
assign q[733]= 16'h32f7;
assign q[734]= 16'h3365;
assign q[735]= 16'h3365;
assign q[736]= 16'h3303;
assign q[737]= 16'h324f;
assign q[738]= 16'h315c;
assign q[739]= 16'h3039;
assign q[740]= 16'h2ef9;
assign q[741]= 16'h2daa;
assign q[742]= 16'h2c5b;
assign q[743]= 16'h2b17;
assign q[744]= 16'h29e6;
assign q[745]= 16'h28ce;
assign q[746]= 16'h27d0;
assign q[747]= 16'h26ea;
assign q[748]= 16'h2617;
assign q[749]= 16'h254e;
assign q[750]= 16'h2484;
assign q[751]= 16'h23ac;
assign q[752]= 16'h22b8;
assign q[753]= 16'h2197;
assign q[754]= 16'h203c;
assign q[755]= 16'h1e96;
assign q[756]= 16'h1c9b;
assign q[757]= 16'h1a3f;
assign q[758]= 16'h177b;
assign q[759]= 16'h144c;
assign q[760]= 16'h10b3;
assign q[761]= 16'hcb5;
assign q[762]= 16'h85b;
assign q[763]= 16'h3b5;
assign q[764]= 16'hfed5;
assign q[765]= 16'hf9d1;
assign q[766]= 16'hf4c2;
assign q[767]= 16'hefc5;
assign q[768]= 16'heaf9;
assign q[769]= 16'he67c;
assign q[770]= 16'he26d;
assign q[771]= 16'hdee9;
assign q[772]= 16'hdc0b;
assign q[773]= 16'hd9ec;
assign q[774]= 16'hd89e;
assign q[775]= 16'hd832;
assign q[776]= 16'hd8af;
assign q[777]= 16'hda1a;
assign q[778]= 16'hdc6f;
assign q[779]= 16'hdfa4;
assign q[780]= 16'he3a9;
assign q[781]= 16'he86a;
assign q[782]= 16'hedcb;
assign q[783]= 16'hf3ad;
assign q[784]= 16'hf9ee;
assign q[785]= 16'h67;
assign q[786]= 16'h6f5;
assign q[787]= 16'hd71;
assign q[788]= 16'h13b4;
assign q[789]= 16'h199f;
assign q[790]= 16'h1f11;
assign q[791]= 16'h23f1;
assign q[792]= 16'h282b;
assign q[793]= 16'h2bb0;
assign q[794]= 16'h2e79;
assign q[795]= 16'h3086;
assign q[796]= 16'h31db;
assign q[797]= 16'h3286;
assign q[798]= 16'h3298;
assign q[799]= 16'h3227;
assign q[800]= 16'h3150;
assign q[801]= 16'h302e;
assign q[802]= 16'h2ee1;
assign q[803]= 16'h2d88;
assign q[804]= 16'h2c3f;
assign q[805]= 16'h2b23;
assign q[806]= 16'h2a49;
assign q[807]= 16'h29c4;
assign q[808]= 16'h29a1;
assign q[809]= 16'h29e4;
assign q[810]= 16'h2a8d;
assign q[811]= 16'h2b95;
assign q[812]= 16'h2ceb;
assign q[813]= 16'h2e7d;
assign q[814]= 16'h302f;
assign q[815]= 16'h31e4;
assign q[816]= 16'h337a;
assign q[817]= 16'h34cf;
assign q[818]= 16'h35bf;
assign q[819]= 16'h3629;
assign q[820]= 16'h35ef;
assign q[821]= 16'h34f7;
assign q[822]= 16'h332e;
assign q[823]= 16'h3087;
assign q[824]= 16'h2cfe;
assign q[825]= 16'h2897;
assign q[826]= 16'h235f;
assign q[827]= 16'h1d6b;
assign q[828]= 16'h16db;
assign q[829]= 16'hfd2;
assign q[830]= 16'h87d;
assign q[831]= 16'h10d;
assign q[832]= 16'hf9b6;
assign q[833]= 16'hf2ad;
assign q[834]= 16'hec28;
assign q[835]= 16'he658;
assign q[836]= 16'he16c;
assign q[837]= 16'hdd8d;
assign q[838]= 16'hdad9;
assign q[839]= 16'hd968;
assign q[840]= 16'hd946;
assign q[841]= 16'hda76;
assign q[842]= 16'hdcec;
assign q[843]= 16'he095;
assign q[844]= 16'he551;
assign q[845]= 16'heaf7;
assign q[846]= 16'hf155;
assign q[847]= 16'hf833;
assign q[848]= 16'hff54;
assign q[849]= 16'h678;
assign q[850]= 16'hd61;
assign q[851]= 16'h13cf;
assign q[852]= 16'h1989;
assign q[853]= 16'h1e5a;
assign q[854]= 16'h2217;
assign q[855]= 16'h249d;
assign q[856]= 16'h25d6;
assign q[857]= 16'h25b6;
assign q[858]= 16'h243e;
assign q[859]= 16'h217c;
assign q[860]= 16'h1d87;
assign q[861]= 16'h1885;
assign q[862]= 16'h12a2;
assign q[863]= 16'hc15;
assign q[864]= 16'h518;
assign q[865]= 16'hfdec;
assign q[866]= 16'hf6d0;
assign q[867]= 16'hf006;
assign q[868]= 16'he9ca;
assign q[869]= 16'he454;
assign q[870]= 16'hdfd6;
assign q[871]= 16'hdc78;
assign q[872]= 16'hda56;
assign q[873]= 16'hd985;
assign q[874]= 16'hda0a;
assign q[875]= 16'hdbe1;
assign q[876]= 16'hdef9;
assign q[877]= 16'he337;
assign q[878]= 16'he877;
assign q[879]= 16'hee8b;
assign q[880]= 16'hf541;
assign q[881]= 16'hfc60;
assign q[882]= 16'h3ae;
assign q[883]= 16'haf2;
assign q[884]= 16'h11f3;
assign q[885]= 16'h187e;
assign q[886]= 16'h1e64;
assign q[887]= 16'h237e;
assign q[888]= 16'h27ae;
assign q[889]= 16'h2ade;
assign q[890]= 16'h2d04;
assign q[891]= 16'h2e1e;
assign q[892]= 16'h2e37;
assign q[893]= 16'h2d61;
assign q[894]= 16'h2bb6;
assign q[895]= 16'h2957;
assign q[896]= 16'h266b;
assign q[897]= 16'h231e;
assign q[898]= 16'h1f9c;
assign q[899]= 16'h1c11;
assign q[900]= 16'h18aa;
assign q[901]= 16'h158d;
assign q[902]= 16'h12de;
assign q[903]= 16'h10b9;
assign q[904]= 16'hf35;
assign q[905]= 16'he60;
assign q[906]= 16'he40;
assign q[907]= 16'hed2;
assign q[908]= 16'h100d;
assign q[909]= 16'h11e0;
assign q[910]= 16'h1433;
assign q[911]= 16'h16eb;
assign q[912]= 16'h19e6;
assign q[913]= 16'h1d03;
assign q[914]= 16'h201e;
assign q[915]= 16'h2315;
assign q[916]= 16'h25c8;
assign q[917]= 16'h2818;
assign q[918]= 16'h29ee;
assign q[919]= 16'h2b38;
assign q[920]= 16'h2be8;
assign q[921]= 16'h2bf9;
assign q[922]= 16'h2b6b;
assign q[923]= 16'h2a47;
assign q[924]= 16'h289b;
assign q[925]= 16'h267a;
assign q[926]= 16'h23fc;
assign q[927]= 16'h213d;
assign q[928]= 16'h1e5c;
assign q[929]= 16'h1b79;
assign q[930]= 16'h18b1;
assign q[931]= 16'h1624;
assign q[932]= 16'h13ec;
assign q[933]= 16'h1221;
assign q[934]= 16'h10d6;
assign q[935]= 16'h1017;
assign q[936]= 16'hfec;
assign q[937]= 16'h1055;
assign q[938]= 16'h114f;
assign q[939]= 16'h12cc;
assign q[940]= 16'h14bd;
assign q[941]= 16'h170c;
assign q[942]= 16'h199e;
assign q[943]= 16'h1c57;
assign q[944]= 16'h1f17;
assign q[945]= 16'h21be;
assign q[946]= 16'h242c;
assign q[947]= 16'h2643;
assign q[948]= 16'h27e6;
assign q[949]= 16'h28fd;
assign q[950]= 16'h2972;
assign q[951]= 16'h2936;
assign q[952]= 16'h283e;
assign q[953]= 16'h2684;
assign q[954]= 16'h240a;
assign q[955]= 16'h20d5;
assign q[956]= 16'h1cef;
assign q[957]= 16'h186a;
assign q[958]= 16'h1359;
assign q[959]= 16'hdd4;
assign q[960]= 16'h7f5;
assign q[961]= 16'h1d7;
assign q[962]= 16'hfb9a;
assign q[963]= 16'hf557;
assign q[964]= 16'hef2c;
assign q[965]= 16'he934;
assign q[966]= 16'he388;
assign q[967]= 16'hde3e;
assign q[968]= 16'hd968;
assign q[969]= 16'hd516;
assign q[970]= 16'hd154;
assign q[971]= 16'hce2b;
assign q[972]= 16'hcb9f;
assign q[973]= 16'hc9b2;
assign q[974]= 16'hc861;
assign q[975]= 16'hc7a8;
assign q[976]= 16'hc781;
assign q[977]= 16'hc7e3;
assign q[978]= 16'hc8c3;
assign q[979]= 16'hca16;
assign q[980]= 16'hcbd0;
assign q[981]= 16'hcde5;
assign q[982]= 16'hd049;
assign q[983]= 16'hd2f1;
assign q[984]= 16'hd5d1;
assign q[985]= 16'hd8e0;
assign q[986]= 16'hdc14;
assign q[987]= 16'hdf64;
assign q[988]= 16'he2c9;
assign q[989]= 16'he63d;
assign q[990]= 16'he9b9;
assign q[991]= 16'hed39;
assign q[992]= 16'hf0b6;
assign q[993]= 16'hf42c;
assign q[994]= 16'hf797;
assign q[995]= 16'hfaf2;
assign q[996]= 16'hfe37;
assign q[997]= 16'h162;
assign q[998]= 16'h46e;
assign q[999]= 16'h756;
assign q[1000]= 16'ha12;
assign q[1001]= 16'hc9c;
assign q[1002]= 16'heef;
assign q[1003]= 16'h1103;
assign q[1004]= 16'h12d2;
assign q[1005]= 16'h1456;
assign q[1006]= 16'h1589;
assign q[1007]= 16'h1666;
assign q[1008]= 16'h16e7;
assign q[1009]= 16'h170a;
assign q[1010]= 16'h16cb;
assign q[1011]= 16'h1629;
assign q[1012]= 16'h1523;
assign q[1013]= 16'h13bb;
assign q[1014]= 16'h11f3;
assign q[1015]= 16'hfcf;
assign q[1016]= 16'hd54;
assign q[1017]= 16'ha88;
assign q[1018]= 16'h775;
assign q[1019]= 16'h424;
assign q[1020]= 16'h9e;
assign q[1021]= 16'hfcf1;
assign q[1022]= 16'hf927;
assign q[1023]= 16'hf54e;
assign q[1024]= 16'hf173;
assign q[1025]= 16'heda5;
assign q[1026]= 16'he9f2;
assign q[1027]= 16'he667;
assign q[1028]= 16'he312;
assign q[1029]= 16'hdfff;
assign q[1030]= 16'hdd3a;
assign q[1031]= 16'hdacd;
assign q[1032]= 16'hd8c4;
assign q[1033]= 16'hd725;
assign q[1034]= 16'hd5f6;
assign q[1035]= 16'hd53d;
assign q[1036]= 16'hd4fd;
assign q[1037]= 16'hd535;
assign q[1038]= 16'hd5e7;
assign q[1039]= 16'hd70e;
assign q[1040]= 16'hd8a6;
assign q[1041]= 16'hdaaa;
assign q[1042]= 16'hdd11;
assign q[1043]= 16'hdfd2;
assign q[1044]= 16'he2e4;
assign q[1045]= 16'he63c;
assign q[1046]= 16'he9ce;
assign q[1047]= 16'hed8e;
assign q[1048]= 16'hf171;
assign q[1049]= 16'hf56b;
assign q[1050]= 16'hf971;
assign q[1051]= 16'hfd78;
assign q[1052]= 16'h175;
assign q[1053]= 16'h563;
assign q[1054]= 16'h938;
assign q[1055]= 16'hcec;
assign q[1056]= 16'h107c;
assign q[1057]= 16'h13e0;
assign q[1058]= 16'h1717;
assign q[1059]= 16'h1a1b;
assign q[1060]= 16'h1cea;
assign q[1061]= 16'h1f82;
assign q[1062]= 16'h21de;
assign q[1063]= 16'h23fd;
assign q[1064]= 16'h25da;
assign q[1065]= 16'h2772;
assign q[1066]= 16'h28c0;
assign q[1067]= 16'h29bf;
assign q[1068]= 16'h2a69;
assign q[1069]= 16'h2ab8;
assign q[1070]= 16'h2aa5;
assign q[1071]= 16'h2a2b;
assign q[1072]= 16'h2941;
assign q[1073]= 16'h27e4;
assign q[1074]= 16'h260e;
assign q[1075]= 16'h23bd;
assign q[1076]= 16'h20ee;
assign q[1077]= 16'h1da4;
assign q[1078]= 16'h19e3;
assign q[1079]= 16'h15b2;
assign q[1080]= 16'h111a;
assign q[1081]= 16'hc2b;
assign q[1082]= 16'h6f5;
assign q[1083]= 16'h18d;
assign q[1084]= 16'hfc0b;
assign q[1085]= 16'hf688;
assign q[1086]= 16'hf120;
assign q[1087]= 16'hebf1;
assign q[1088]= 16'he71a;
assign q[1089]= 16'he2b8;
assign q[1090]= 16'hdee7;
assign q[1091]= 16'hdbc3;
assign q[1092]= 16'hd962;
assign q[1093]= 16'hd7d7;
assign q[1094]= 16'hd732;
assign q[1095]= 16'hd77c;
assign q[1096]= 16'hd8b8;
assign q[1097]= 16'hdae2;
assign q[1098]= 16'hddf1;
assign q[1099]= 16'he1d5;
assign q[1100]= 16'he679;
assign q[1101]= 16'hebbf;
assign q[1102]= 16'hf189;
assign q[1103]= 16'hf7b1;
assign q[1104]= 16'hfe11;
assign q[1105]= 16'h47e;
assign q[1106]= 16'had2;
assign q[1107]= 16'h10e2;
assign q[1108]= 16'h168b;
assign q[1109]= 16'h1ba8;
assign q[1110]= 16'h201e;
assign q[1111]= 16'h23d3;
assign q[1112]= 16'h26b8;
assign q[1113]= 16'h28c2;
assign q[1114]= 16'h29f0;
assign q[1115]= 16'h2a45;
assign q[1116]= 16'h29d0;
assign q[1117]= 16'h28a2;
assign q[1118]= 16'h26d6;
assign q[1119]= 16'h248a;
assign q[1120]= 16'h21e1;
assign q[1121]= 16'h1eff;
assign q[1122]= 16'h1c0a;
assign q[1123]= 16'h1929;
assign q[1124]= 16'h167f;
assign q[1125]= 16'h142d;
assign q[1126]= 16'h124e;
assign q[1127]= 16'h10fa;
assign q[1128]= 16'h103f;
assign q[1129]= 16'h1027;
assign q[1130]= 16'h10b3;
assign q[1131]= 16'h11dd;
assign q[1132]= 16'h1396;
assign q[1133]= 16'h15ca;
assign q[1134]= 16'h185f;
assign q[1135]= 16'h1b35;
assign q[1136]= 16'h1e29;
assign q[1137]= 16'h2115;
assign q[1138]= 16'h23d3;
assign q[1139]= 16'h263d;
assign q[1140]= 16'h2830;
assign q[1141]= 16'h298b;
assign q[1142]= 16'h2a33;
assign q[1143]= 16'h2a13;
assign q[1144]= 16'h291d;
assign q[1145]= 16'h2748;
assign q[1146]= 16'h2495;
assign q[1147]= 16'h210b;
assign q[1148]= 16'h1cbb;
assign q[1149]= 16'h17b9;
assign q[1150]= 16'h1222;
assign q[1151]= 16'hc17;
assign q[1152]= 16'h5bb;
assign q[1153]= 16'hff37;
assign q[1154]= 16'hf8b1;
assign q[1155]= 16'hf251;
assign q[1156]= 16'hec3e;
assign q[1157]= 16'he69a;
assign q[1158]= 16'he186;
assign q[1159]= 16'hdd19;
assign q[1160]= 16'hd96a;
assign q[1161]= 16'hd686;
assign q[1162]= 16'hd474;
assign q[1163]= 16'hd335;
assign q[1164]= 16'hd2c5;
assign q[1165]= 16'hd319;
assign q[1166]= 16'hd420;
assign q[1167]= 16'hd5c6;
assign q[1168]= 16'hd7f3;
assign q[1169]= 16'hda8d;
assign q[1170]= 16'hdd78;
assign q[1171]= 16'he098;
assign q[1172]= 16'he3d1;
assign q[1173]= 16'he70a;
assign q[1174]= 16'hea2a;
assign q[1175]= 16'hed1d;
assign q[1176]= 16'hefd0;
assign q[1177]= 16'hf237;
assign q[1178]= 16'hf445;
assign q[1179]= 16'hf5f6;
assign q[1180]= 16'hf745;
assign q[1181]= 16'hf832;
assign q[1182]= 16'hf8c0;
assign q[1183]= 16'hf8f3;
assign q[1184]= 16'hf8d4;
assign q[1185]= 16'hf868;
assign q[1186]= 16'hf7ba;
assign q[1187]= 16'hf6d2;
assign q[1188]= 16'hf5b8;
assign q[1189]= 16'hf474;
assign q[1190]= 16'hf30e;
assign q[1191]= 16'hf18d;
assign q[1192]= 16'heff5;
assign q[1193]= 16'hee4b;
assign q[1194]= 16'hec93;
assign q[1195]= 16'head0;
assign q[1196]= 16'he905;
assign q[1197]= 16'he733;
assign q[1198]= 16'he55e;
assign q[1199]= 16'he387;
assign q[1200]= 16'he1b1;
assign q[1201]= 16'hdfe1;
assign q[1202]= 16'hde1a;
assign q[1203]= 16'hdc60;
assign q[1204]= 16'hdab8;
assign q[1205]= 16'hd928;
assign q[1206]= 16'hd7b5;
assign q[1207]= 16'hd663;
assign q[1208]= 16'hd539;
assign q[1209]= 16'hd438;
assign q[1210]= 16'hd366;
assign q[1211]= 16'hd2c3;
assign q[1212]= 16'hd250;
assign q[1213]= 16'hd20d;
assign q[1214]= 16'hd1f6;
assign q[1215]= 16'hd209;
assign q[1216]= 16'hd240;
assign q[1217]= 16'hd294;
assign q[1218]= 16'hd301;
assign q[1219]= 16'hd37e;
assign q[1220]= 16'hd405;
assign q[1221]= 16'hd48f;
assign q[1222]= 16'hd517;
assign q[1223]= 16'hd59a;
assign q[1224]= 16'hd616;
assign q[1225]= 16'hd68a;
assign q[1226]= 16'hd6f9;
assign q[1227]= 16'hd768;
assign q[1228]= 16'hd7de;
assign q[1229]= 16'hd864;
assign q[1230]= 16'hd906;
assign q[1231]= 16'hd9cf;
assign q[1232]= 16'hdacd;
assign q[1233]= 16'hdc0d;
assign q[1234]= 16'hdd9c;
assign q[1235]= 16'hdf85;
assign q[1236]= 16'he1d3;
assign q[1237]= 16'he48c;
assign q[1238]= 16'he7b4;
assign q[1239]= 16'heb4a;
assign q[1240]= 16'hef4a;
assign q[1241]= 16'hf3ac;
assign q[1242]= 16'hf862;
assign q[1243]= 16'hfd5b;
assign q[1244]= 16'h280;
assign q[1245]= 16'h7b9;
assign q[1246]= 16'hceb;
assign q[1247]= 16'h11f8;
assign q[1248]= 16'h16c0;
assign q[1249]= 16'h1b25;
assign q[1250]= 16'h1f09;
assign q[1251]= 16'h224f;
assign q[1252]= 16'h24e0;
assign q[1253]= 16'h26a7;
assign q[1254]= 16'h2794;
assign q[1255]= 16'h279c;
assign q[1256]= 16'h26bc;
assign q[1257]= 16'h24f4;
assign q[1258]= 16'h224c;
assign q[1259]= 16'h1ed4;
assign q[1260]= 16'h1a9e;
assign q[1261]= 16'h15c4;
assign q[1262]= 16'h1062;
assign q[1263]= 16'ha99;
assign q[1264]= 16'h48c;
assign q[1265]= 16'hfe60;
assign q[1266]= 16'hf839;
assign q[1267]= 16'hf23a;
assign q[1268]= 16'hec84;
assign q[1269]= 16'he738;
assign q[1270]= 16'he26e;
assign q[1271]= 16'hde3f;
assign q[1272]= 16'hdabb;
assign q[1273]= 16'hd7ef;
assign q[1274]= 16'hd5e0;
assign q[1275]= 16'hd490;
assign q[1276]= 16'hd3fc;
assign q[1277]= 16'hd41a;
assign q[1278]= 16'hd4de;
assign q[1279]= 16'hd636;
assign q[1280]= 16'hd80f;
assign q[1281]= 16'hda54;
assign q[1282]= 16'hdced;
assign q[1283]= 16'hdfc3;
assign q[1284]= 16'he2be;
assign q[1285]= 16'he5c7;
assign q[1286]= 16'he8ca;
assign q[1287]= 16'hebb3;
assign q[1288]= 16'hee70;
assign q[1289]= 16'hf0f4;
assign q[1290]= 16'hf333;
assign q[1291]= 16'hf522;
assign q[1292]= 16'hf6bd;
assign q[1293]= 16'hf7fe;
assign q[1294]= 16'hf8e4;
assign q[1295]= 16'hf971;
assign q[1296]= 16'hf9a6;
assign q[1297]= 16'hf988;
assign q[1298]= 16'hf91d;
assign q[1299]= 16'hf86b;
assign q[1300]= 16'hf77b;
assign q[1301]= 16'hf656;
assign q[1302]= 16'hf505;
assign q[1303]= 16'hf393;
assign q[1304]= 16'hf20a;
assign q[1305]= 16'hf076;
assign q[1306]= 16'heee4;
assign q[1307]= 16'hed5e;
assign q[1308]= 16'hebf2;
assign q[1309]= 16'heaad;
assign q[1310]= 16'he999;
assign q[1311]= 16'he8c5;
assign q[1312]= 16'he83c;
assign q[1313]= 16'he809;
assign q[1314]= 16'he836;
assign q[1315]= 16'he8cb;
assign q[1316]= 16'he9cf;
assign q[1317]= 16'heb46;
assign q[1318]= 16'hed33;
assign q[1319]= 16'hef94;
assign q[1320]= 16'hf267;
assign q[1321]= 16'hf5a2;
assign q[1322]= 16'hf93d;
assign q[1323]= 16'hfd29;
assign q[1324]= 16'h154;
assign q[1325]= 16'h5ae;
assign q[1326]= 16'ha1f;
assign q[1327]= 16'he8f;
assign q[1328]= 16'h12e6;
assign q[1329]= 16'h170b;
assign q[1330]= 16'h1ae3;
assign q[1331]= 16'h1e58;
assign q[1332]= 16'h2152;
assign q[1333]= 16'h23be;
assign q[1334]= 16'h258c;
assign q[1335]= 16'h26af;
assign q[1336]= 16'h271f;
assign q[1337]= 16'h26d8;
assign q[1338]= 16'h25dd;
assign q[1339]= 16'h2434;
assign q[1340]= 16'h21e8;
assign q[1341]= 16'h1f09;
assign q[1342]= 16'h1bab;
assign q[1343]= 16'h17e5;
assign q[1344]= 16'h13d1;
assign q[1345]= 16'hf8a;
assign q[1346]= 16'hb2d;
assign q[1347]= 16'h6d6;
assign q[1348]= 16'h29e;
assign q[1349]= 16'hfea1;
assign q[1350]= 16'hfaf1;
assign q[1351]= 16'hf7a3;
assign q[1352]= 16'hf4c4;
assign q[1353]= 16'hf25d;
assign q[1354]= 16'hf074;
assign q[1355]= 16'hef08;
assign q[1356]= 16'hee14;
assign q[1357]= 16'hed90;
assign q[1358]= 16'hed6c;
assign q[1359]= 16'hed9a;
assign q[1360]= 16'hee06;
assign q[1361]= 16'hee9c;
assign q[1362]= 16'hef45;
assign q[1363]= 16'hefed;
assign q[1364]= 16'hf07e;
assign q[1365]= 16'hf0e7;
assign q[1366]= 16'hf117;
assign q[1367]= 16'hf101;
assign q[1368]= 16'hf09c;
assign q[1369]= 16'hefe3;
assign q[1370]= 16'heed3;
assign q[1371]= 16'hed71;
assign q[1372]= 16'hebc3;
assign q[1373]= 16'he9d4;
assign q[1374]= 16'he7b2;
assign q[1375]= 16'he56d;
assign q[1376]= 16'he319;
assign q[1377]= 16'he0c9;
assign q[1378]= 16'hde92;
assign q[1379]= 16'hdc89;
assign q[1380]= 16'hdac2;
assign q[1381]= 16'hd94e;
assign q[1382]= 16'hd83f;
assign q[1383]= 16'hd7a1;
assign q[1384]= 16'hd780;
assign q[1385]= 16'hd7e3;
assign q[1386]= 16'hd8ce;
assign q[1387]= 16'hda40;
assign q[1388]= 16'hdc38;
assign q[1389]= 16'hdeae;
assign q[1390]= 16'he19a;
assign q[1391]= 16'he4ee;
assign q[1392]= 16'he89e;
assign q[1393]= 16'hec98;
assign q[1394]= 16'hf0cb;
assign q[1395]= 16'hf523;
assign q[1396]= 16'hf98e;
assign q[1397]= 16'hfdf9;
assign q[1398]= 16'h24e;
assign q[1399]= 16'h67e;
assign q[1400]= 16'ha75;
assign q[1401]= 16'he24;
assign q[1402]= 16'h117b;
assign q[1403]= 16'h146d;
assign q[1404]= 16'h16ef;
assign q[1405]= 16'h18f6;
assign q[1406]= 16'h1a7c;
assign q[1407]= 16'h1b7a;
assign q[1408]= 16'h1bec;
assign q[1409]= 16'h1bd1;
assign q[1410]= 16'h1b2a;
assign q[1411]= 16'h19f8;
assign q[1412]= 16'h1841;
assign q[1413]= 16'h160a;
assign q[1414]= 16'h135e;
assign q[1415]= 16'h1045;
assign q[1416]= 16'hccd;
assign q[1417]= 16'h904;
assign q[1418]= 16'h4f9;
assign q[1419]= 16'hbf;
assign q[1420]= 16'hfc69;
assign q[1421]= 16'hf809;
assign q[1422]= 16'hf3b4;
assign q[1423]= 16'hef7f;
assign q[1424]= 16'heb7f;
assign q[1425]= 16'he7c9;
assign q[1426]= 16'he471;
assign q[1427]= 16'he189;
assign q[1428]= 16'hdf24;
assign q[1429]= 16'hdd50;
assign q[1430]= 16'hdc1a;
assign q[1431]= 16'hdb8d;
assign q[1432]= 16'hdbb1;
assign q[1433]= 16'hdc8a;
assign q[1434]= 16'hde19;
assign q[1435]= 16'he05b;
assign q[1436]= 16'he34c;
assign q[1437]= 16'he6e3;
assign q[1438]= 16'heb12;
assign q[1439]= 16'hefcc;
assign q[1440]= 16'hf4fd;
assign q[1441]= 16'hfa93;
assign q[1442]= 16'h77;
assign q[1443]= 16'h691;
assign q[1444]= 16'hcc9;
assign q[1445]= 16'h1306;
assign q[1446]= 16'h192e;
assign q[1447]= 16'h1f26;
assign q[1448]= 16'h24d8;
assign q[1449]= 16'h2a2c;
assign q[1450]= 16'h2f0a;
assign q[1451]= 16'h3361;
assign q[1452]= 16'h371d;
assign q[1453]= 16'h3a2f;
assign q[1454]= 16'h3c8a;
assign q[1455]= 16'h3e24;
assign q[1456]= 16'h3ef6;
assign q[1457]= 16'h3efc;
assign q[1458]= 16'h3e36;
assign q[1459]= 16'h3ca5;
assign q[1460]= 16'h3a4f;
assign q[1461]= 16'h373c;
assign q[1462]= 16'h3378;
assign q[1463]= 16'h2f11;
assign q[1464]= 16'h2a19;
assign q[1465]= 16'h24a4;
assign q[1466]= 16'h1ec8;
assign q[1467]= 16'h189e;
assign q[1468]= 16'h123f;
assign q[1469]= 16'hbc7;
assign q[1470]= 16'h554;
assign q[1471]= 16'hff02;
assign q[1472]= 16'hf8ee;
assign q[1473]= 16'hf334;
assign q[1474]= 16'hedf1;
assign q[1475]= 16'he93f;
assign q[1476]= 16'he534;
assign q[1477]= 16'he1e7;
assign q[1478]= 16'hdf68;
assign q[1479]= 16'hddc5;
assign q[1480]= 16'hdd07;
assign q[1481]= 16'hdd34;
assign q[1482]= 16'hde4b;
assign q[1483]= 16'he047;
assign q[1484]= 16'he31e;
assign q[1485]= 16'he6c2;
assign q[1486]= 16'heb1f;
assign q[1487]= 16'hf01e;
assign q[1488]= 16'hf5a5;
assign q[1489]= 16'hfb95;
assign q[1490]= 16'h1cf;
assign q[1491]= 16'h831;
assign q[1492]= 16'he9b;
assign q[1493]= 16'h14eb;
assign q[1494]= 16'h1b01;
assign q[1495]= 16'h20bf;
assign q[1496]= 16'h260c;
assign q[1497]= 16'h2acf;
assign q[1498]= 16'h2ef6;
assign q[1499]= 16'h3274;
assign q[1500]= 16'h353e;
assign q[1501]= 16'h374f;
assign q[1502]= 16'h38aa;
assign q[1503]= 16'h3952;
assign q[1504]= 16'h3950;
assign q[1505]= 16'h38b2;
assign q[1506]= 16'h3788;
assign q[1507]= 16'h35e2;
assign q[1508]= 16'h33d4;
assign q[1509]= 16'h3172;
assign q[1510]= 16'h2ed0;
assign q[1511]= 16'h2bff;
assign q[1512]= 16'h2910;
assign q[1513]= 16'h2611;
assign q[1514]= 16'h230e;
assign q[1515]= 16'h200e;
assign q[1516]= 16'h1d16;
assign q[1517]= 16'h1a29;
assign q[1518]= 16'h1744;
assign q[1519]= 16'h1464;
assign q[1520]= 16'h1183;
assign q[1521]= 16'he99;
assign q[1522]= 16'hb9e;
assign q[1523]= 16'h88a;
assign q[1524]= 16'h556;
assign q[1525]= 16'h1fb;
assign q[1526]= 16'hfe78;
assign q[1527]= 16'hfac8;
assign q[1528]= 16'hf6f1;
assign q[1529]= 16'hf2f7;
assign q[1530]= 16'heee5;
assign q[1531]= 16'heac8;
assign q[1532]= 16'he6b0;
assign q[1533]= 16'he2b2;
assign q[1534]= 16'hdee4;
assign q[1535]= 16'hdb5c;
assign q[1536]= 16'hd835;
assign q[1537]= 16'hd586;
assign q[1538]= 16'hd367;
assign q[1539]= 16'hd1ec;
assign q[1540]= 16'hd128;
assign q[1541]= 16'hd129;
assign q[1542]= 16'hd1f8;
assign q[1543]= 16'hd39a;
assign q[1544]= 16'hd60f;
assign q[1545]= 16'hd94e;
assign q[1546]= 16'hdd4b;
assign q[1547]= 16'he1f4;
assign q[1548]= 16'he732;
assign q[1549]= 16'hecea;
assign q[1550]= 16'hf2fb;
assign q[1551]= 16'hf945;
assign q[1552]= 16'hffa4;
assign q[1553]= 16'h5f3;
assign q[1554]= 16'hc12;
assign q[1555]= 16'h11dd;
assign q[1556]= 16'h1737;
assign q[1557]= 16'h1c06;
assign q[1558]= 16'h2033;
assign q[1559]= 16'h23ad;
assign q[1560]= 16'h266b;
assign q[1561]= 16'h2865;
assign q[1562]= 16'h299e;
assign q[1563]= 16'h2a1c;
assign q[1564]= 16'h29e9;
assign q[1565]= 16'h2917;
assign q[1566]= 16'h27b8;
assign q[1567]= 16'h25e5;
assign q[1568]= 16'h23b7;
assign q[1569]= 16'h2147;
assign q[1570]= 16'h1eb0;
assign q[1571]= 16'h1c0c;
assign q[1572]= 16'h1972;
assign q[1573]= 16'h16f7;
assign q[1574]= 16'h14ae;
assign q[1575]= 16'h12a6;
assign q[1576]= 16'h10e8;
assign q[1577]= 16'hf7b;
assign q[1578]= 16'he61;
assign q[1579]= 16'hd99;
assign q[1580]= 16'hd1c;
assign q[1581]= 16'hce3;
assign q[1582]= 16'hce1;
assign q[1583]= 16'hd09;
assign q[1584]= 16'hd4c;
assign q[1585]= 16'hd9a;
assign q[1586]= 16'hde3;
assign q[1587]= 16'he17;
assign q[1588]= 16'he26;
assign q[1589]= 16'he05;
assign q[1590]= 16'hda6;
assign q[1591]= 16'hd00;
assign q[1592]= 16'hc0c;
assign q[1593]= 16'hac5;
assign q[1594]= 16'h927;
assign q[1595]= 16'h732;
assign q[1596]= 16'h4e7;
assign q[1597]= 16'h24a;
assign q[1598]= 16'hff60;
assign q[1599]= 16'hfc2f;
assign q[1600]= 16'hf8be;
assign q[1601]= 16'hf517;
assign q[1602]= 16'hf144;
assign q[1603]= 16'hed4f;
assign q[1604]= 16'he942;
assign q[1605]= 16'he52b;
assign q[1606]= 16'he116;
assign q[1607]= 16'hdd0e;
assign q[1608]= 16'hd923;
assign q[1609]= 16'hd562;
assign q[1610]= 16'hd1da;
assign q[1611]= 16'hce99;
assign q[1612]= 16'hcbae;
assign q[1613]= 16'hc929;
assign q[1614]= 16'hc718;
assign q[1615]= 16'hc58b;
assign q[1616]= 16'hc48e;
assign q[1617]= 16'hc42d;
assign q[1618]= 16'hc474;
assign q[1619]= 16'hc56b;
assign q[1620]= 16'hc716;
assign q[1621]= 16'hc978;
assign q[1622]= 16'hcc91;
assign q[1623]= 16'hd05a;
assign q[1624]= 16'hd4ca;
assign q[1625]= 16'hd9d4;
assign q[1626]= 16'hdf65;
assign q[1627]= 16'he568;
assign q[1628]= 16'hebc2;
assign q[1629]= 16'hf256;
assign q[1630]= 16'hf904;
assign q[1631]= 16'hffab;
assign q[1632]= 16'h625;
assign q[1633]= 16'hc53;
assign q[1634]= 16'h1212;
assign q[1635]= 16'h1741;
assign q[1636]= 16'h1bc4;
assign q[1637]= 16'h1f82;
assign q[1638]= 16'h2267;
assign q[1639]= 16'h2466;
assign q[1640]= 16'h2577;
assign q[1641]= 16'h2599;
assign q[1642]= 16'h24d2;
assign q[1643]= 16'h2330;
assign q[1644]= 16'h20c5;
assign q[1645]= 16'h1dac;
assign q[1646]= 16'h1a03;
assign q[1647]= 16'h15ed;
assign q[1648]= 16'h1191;
assign q[1649]= 16'hd16;
assign q[1650]= 16'h8a5;
assign q[1651]= 16'h466;
assign q[1652]= 16'h80;
assign q[1653]= 16'hfd15;
assign q[1654]= 16'hfa43;
assign q[1655]= 16'hf823;
assign q[1656]= 16'hf6c8;
assign q[1657]= 16'hf63c;
assign q[1658]= 16'hf686;
assign q[1659]= 16'hf7a3;
assign q[1660]= 16'hf988;
assign q[1661]= 16'hfc26;
assign q[1662]= 16'hff67;
assign q[1663]= 16'h32f;
assign q[1664]= 16'h760;
assign q[1665]= 16'hbd9;
assign q[1666]= 16'h1075;
assign q[1667]= 16'h1512;
assign q[1668]= 16'h198c;
assign q[1669]= 16'h1dc1;
assign q[1670]= 16'h2196;
assign q[1671]= 16'h24f0;
assign q[1672]= 16'h27ba;
assign q[1673]= 16'h29e5;
assign q[1674]= 16'h2b66;
assign q[1675]= 16'h2c3b;
assign q[1676]= 16'h2c64;
assign q[1677]= 16'h2be8;
assign q[1678]= 16'h2ad2;
assign q[1679]= 16'h2934;
assign q[1680]= 16'h271f;
assign q[1681]= 16'h24a9;
assign q[1682]= 16'h21eb;
assign q[1683]= 16'h1efc;
assign q[1684]= 16'h1bf4;
assign q[1685]= 16'h18eb;
assign q[1686]= 16'h15f5;
assign q[1687]= 16'h1327;
assign q[1688]= 16'h1091;
assign q[1689]= 16'he40;
assign q[1690]= 16'hc3f;
assign q[1691]= 16'ha94;
assign q[1692]= 16'h944;
assign q[1693]= 16'h84f;
assign q[1694]= 16'h7b4;
assign q[1695]= 16'h76d;
assign q[1696]= 16'h776;
assign q[1697]= 16'h7c5;
assign q[1698]= 16'h853;
assign q[1699]= 16'h916;
assign q[1700]= 16'ha03;
assign q[1701]= 16'hb11;
assign q[1702]= 16'hc36;
assign q[1703]= 16'hd69;
assign q[1704]= 16'hea0;
assign q[1705]= 16'hfd4;
assign q[1706]= 16'h10fb;
assign q[1707]= 16'h1210;
assign q[1708]= 16'h1309;
assign q[1709]= 16'h13e1;
assign q[1710]= 16'h1491;
assign q[1711]= 16'h1513;
assign q[1712]= 16'h1561;
assign q[1713]= 16'h1575;
assign q[1714]= 16'h154b;
assign q[1715]= 16'h14dd;
assign q[1716]= 16'h1428;
assign q[1717]= 16'h132a;
assign q[1718]= 16'h11e1;
assign q[1719]= 16'h104f;
assign q[1720]= 16'he76;
assign q[1721]= 16'hc5b;
assign q[1722]= 16'ha06;
assign q[1723]= 16'h780;
assign q[1724]= 16'h4d7;
assign q[1725]= 16'h218;
assign q[1726]= 16'hff56;
assign q[1727]= 16'hfca3;
assign q[1728]= 16'hfa13;
assign q[1729]= 16'hf7bb;
assign q[1730]= 16'hf5b2;
assign q[1731]= 16'hf40b;
assign q[1732]= 16'hf2da;
assign q[1733]= 16'hf22f;
assign q[1734]= 16'hf219;
assign q[1735]= 16'hf2a1;
assign q[1736]= 16'hf3cd;
assign q[1737]= 16'hf59e;
assign q[1738]= 16'hf80d;
assign q[1739]= 16'hfb11;
assign q[1740]= 16'hfe9b;
assign q[1741]= 16'h293;
assign q[1742]= 16'h6e2;
assign q[1743]= 16'hb6a;
assign q[1744]= 16'h1008;
assign q[1745]= 16'h149b;
assign q[1746]= 16'h18fe;
assign q[1747]= 16'h1d0d;
assign q[1748]= 16'h20a7;
assign q[1749]= 16'h23ac;
assign q[1750]= 16'h2601;
assign q[1751]= 16'h2791;
assign q[1752]= 16'h284d;
assign q[1753]= 16'h282b;
assign q[1754]= 16'h272b;
assign q[1755]= 16'h2553;
assign q[1756]= 16'h22b2;
assign q[1757]= 16'h1f5c;
assign q[1758]= 16'h1b6e;
assign q[1759]= 16'h1708;
assign q[1760]= 16'h1250;
assign q[1761]= 16'hd6e;
assign q[1762]= 16'h88d;
assign q[1763]= 16'h3d7;
assign q[1764]= 16'hff74;
assign q[1765]= 16'hfb87;
assign q[1766]= 16'hf832;
assign q[1767]= 16'hf58e;
assign q[1768]= 16'hf3af;
assign q[1769]= 16'hf29f;
assign q[1770]= 16'hf262;
assign q[1771]= 16'hf2f0;
assign q[1772]= 16'hf43c;
assign q[1773]= 16'hf62f;
assign q[1774]= 16'hf8ad;
assign q[1775]= 16'hfb92;
assign q[1776]= 16'hfeb8;
assign q[1777]= 16'h1f2;
assign q[1778]= 16'h517;
assign q[1779]= 16'h7fd;
assign q[1780]= 16'ha79;
assign q[1781]= 16'hc68;
assign q[1782]= 16'hdab;
assign q[1783]= 16'he2b;
assign q[1784]= 16'hdd6;
assign q[1785]= 16'hca7;
assign q[1786]= 16'ha9e;
assign q[1787]= 16'h7c7;
assign q[1788]= 16'h435;
assign q[1789]= 16'h4;
assign q[1790]= 16'hfb56;
assign q[1791]= 16'hf654;
assign q[1792]= 16'hf128;
assign q[1793]= 16'hec03;
assign q[1794]= 16'he713;
assign q[1795]= 16'he286;
assign q[1796]= 16'hde87;
assign q[1797]= 16'hdb3a;
assign q[1798]= 16'hd8c0;
assign q[1799]= 16'hd72f;
assign q[1800]= 16'hd697;
assign q[1801]= 16'hd6fd;
assign q[1802]= 16'hd85d;
assign q[1803]= 16'hdaaa;
assign q[1804]= 16'hddce;
assign q[1805]= 16'he1aa;
assign q[1806]= 16'he618;
assign q[1807]= 16'heaef;
assign q[1808]= 16'heffe;
assign q[1809]= 16'hf515;
assign q[1810]= 16'hfa03;
assign q[1811]= 16'hfe98;
assign q[1812]= 16'h2a8;
assign q[1813]= 16'h60d;
assign q[1814]= 16'h8a6;
assign q[1815]= 16'ha5b;
assign q[1816]= 16'hb1d;
assign q[1817]= 16'hae4;
assign q[1818]= 16'h9b4;
assign q[1819]= 16'h799;
assign q[1820]= 16'h4a8;
assign q[1821]= 16'h100;
assign q[1822]= 16'hfcc5;
assign q[1823]= 16'hf81f;
assign q[1824]= 16'hf33e;
assign q[1825]= 16'hee50;
assign q[1826]= 16'he987;
assign q[1827]= 16'he512;
assign q[1828]= 16'he11d;
assign q[1829]= 16'hddd2;
assign q[1830]= 16'hdb52;
assign q[1831]= 16'hd9b8;
assign q[1832]= 16'hd919;
assign q[1833]= 16'hd97f;
assign q[1834]= 16'hdaee;
assign q[1835]= 16'hdd60;
assign q[1836]= 16'he0c8;
assign q[1837]= 16'he510;
assign q[1838]= 16'hea1e;
assign q[1839]= 16'hefcf;
assign q[1840]= 16'hf601;
assign q[1841]= 16'hfc8a;
assign q[1842]= 16'h340;
assign q[1843]= 16'h9ff;
assign q[1844]= 16'h109c;
assign q[1845]= 16'h16f4;
assign q[1846]= 16'h1ce6;
assign q[1847]= 16'h2256;
assign q[1848]= 16'h272d;
assign q[1849]= 16'h2b5d;
assign q[1850]= 16'h2ed9;
assign q[1851]= 16'h319e;
assign q[1852]= 16'h33ae;
assign q[1853]= 16'h350f;
assign q[1854]= 16'h35cf;
assign q[1855]= 16'h35fe;
assign q[1856]= 16'h35ae;
assign q[1857]= 16'h34f6;
assign q[1858]= 16'h33ec;
assign q[1859]= 16'h32a9;
assign q[1860]= 16'h3143;
assign q[1861]= 16'h2fd0;
assign q[1862]= 16'h2e63;
assign q[1863]= 16'h2d0e;
assign q[1864]= 16'h2bde;
assign q[1865]= 16'h2add;
assign q[1866]= 16'h2a13;
assign q[1867]= 16'h2983;
assign q[1868]= 16'h292c;
assign q[1869]= 16'h290d;
assign q[1870]= 16'h291f;
assign q[1871]= 16'h295a;
assign q[1872]= 16'h29b5;
assign q[1873]= 16'h2a24;
assign q[1874]= 16'h2a9d;
assign q[1875]= 16'h2b13;
assign q[1876]= 16'h2b7c;
assign q[1877]= 16'h2bcc;
assign q[1878]= 16'h2bfa;
assign q[1879]= 16'h2bfe;
assign q[1880]= 16'h2bd2;
assign q[1881]= 16'h2b6f;
assign q[1882]= 16'h2ad5;
assign q[1883]= 16'h29ff;
assign q[1884]= 16'h28f0;
assign q[1885]= 16'h27a8;
assign q[1886]= 16'h2629;
assign q[1887]= 16'h2478;
assign q[1888]= 16'h229a;
assign q[1889]= 16'h2092;
assign q[1890]= 16'h1e67;
assign q[1891]= 16'h1c1e;
assign q[1892]= 16'h19bd;
assign q[1893]= 16'h1749;
assign q[1894]= 16'h14c8;
assign q[1895]= 16'h1240;
assign q[1896]= 16'hfb6;
assign q[1897]= 16'hd2d;
assign q[1898]= 16'haac;
assign q[1899]= 16'h837;
assign q[1900]= 16'h5d1;
assign q[1901]= 16'h37f;
assign q[1902]= 16'h146;
assign q[1903]= 16'hff2a;
assign q[1904]= 16'hfd2c;
assign q[1905]= 16'hfb52;
assign q[1906]= 16'hf99f;
assign q[1907]= 16'hf815;
assign q[1908]= 16'hf6b7;
assign q[1909]= 16'hf587;
assign q[1910]= 16'hf485;
assign q[1911]= 16'hf3b1;
assign q[1912]= 16'hf30b;
assign q[1913]= 16'hf291;
assign q[1914]= 16'hf23f;
assign q[1915]= 16'hf211;
assign q[1916]= 16'hf203;
assign q[1917]= 16'hf20d;
assign q[1918]= 16'hf229;
assign q[1919]= 16'hf24e;
assign q[1920]= 16'hf276;
assign q[1921]= 16'hf296;
assign q[1922]= 16'hf2a6;
assign q[1923]= 16'hf29f;
assign q[1924]= 16'hf278;
assign q[1925]= 16'hf22a;
assign q[1926]= 16'hf1b1;
assign q[1927]= 16'hf106;
assign q[1928]= 16'hf029;
assign q[1929]= 16'hef17;
assign q[1930]= 16'hedd2;
assign q[1931]= 16'hec5c;
assign q[1932]= 16'heab9;
assign q[1933]= 16'he8f1;
assign q[1934]= 16'he70a;
assign q[1935]= 16'he50f;
assign q[1936]= 16'he309;
assign q[1937]= 16'he103;
assign q[1938]= 16'hdf0a;
assign q[1939]= 16'hdd29;
assign q[1940]= 16'hdb6c;
assign q[1941]= 16'hd9dd;
assign q[1942]= 16'hd888;
assign q[1943]= 16'hd775;
assign q[1944]= 16'hd6ac;
assign q[1945]= 16'hd633;
assign q[1946]= 16'hd60d;
assign q[1947]= 16'hd63f;
assign q[1948]= 16'hd6c7;
assign q[1949]= 16'hd7a5;
assign q[1950]= 16'hd8d5;
assign q[1951]= 16'hda53;
assign q[1952]= 16'hdc19;
assign q[1953]= 16'hde1e;
assign q[1954]= 16'he05a;
assign q[1955]= 16'he2c4;
assign q[1956]= 16'he553;
assign q[1957]= 16'he7fc;
assign q[1958]= 16'heab5;
assign q[1959]= 16'hed76;
assign q[1960]= 16'hf035;
assign q[1961]= 16'hf2ea;
assign q[1962]= 16'hf58e;
assign q[1963]= 16'hf81a;
assign q[1964]= 16'hfa8a;
assign q[1965]= 16'hfcd8;
assign q[1966]= 16'hff02;
assign q[1967]= 16'h105;
assign q[1968]= 16'h2e1;
assign q[1969]= 16'h495;
assign q[1970]= 16'h621;
assign q[1971]= 16'h787;
assign q[1972]= 16'h8c8;
assign q[1973]= 16'h9e5;
assign q[1974]= 16'hae2;
assign q[1975]= 16'hbbf;
assign q[1976]= 16'hc80;
assign q[1977]= 16'hd27;
assign q[1978]= 16'hdb6;
assign q[1979]= 16'he2f;
assign q[1980]= 16'he94;
assign q[1981]= 16'hee7;
assign q[1982]= 16'hf29;
assign q[1983]= 16'hf5d;
assign q[1984]= 16'hf82;
assign q[1985]= 16'hf9b;
assign q[1986]= 16'hfaa;
assign q[1987]= 16'hfae;
assign q[1988]= 16'hfaa;
assign q[1989]= 16'hf9e;
assign q[1990]= 16'hf8c;
assign q[1991]= 16'hf75;
assign q[1992]= 16'hf5a;
assign q[1993]= 16'hf3d;
assign q[1994]= 16'hf1e;
assign q[1995]= 16'hf00;
assign q[1996]= 16'hee3;
assign q[1997]= 16'hec7;
assign q[1998]= 16'heae;
assign q[1999]= 16'he98;
assign q[2000]= 16'he86;
assign q[2001]= 16'he78;
assign q[2002]= 16'he6d;
assign q[2003]= 16'he66;
assign q[2004]= 16'he61;
assign q[2005]= 16'he5f;
assign q[2006]= 16'he5e;
assign q[2007]= 16'he5e;
assign q[2008]= 16'he5d;
assign q[2009]= 16'he5c;
assign q[2010]= 16'he59;
assign q[2011]= 16'he55;
assign q[2012]= 16'he50;
assign q[2013]= 16'he49;
assign q[2014]= 16'he42;
assign q[2015]= 16'he3d;
assign q[2016]= 16'he3b;
assign q[2017]= 16'he3e;
assign q[2018]= 16'he49;
assign q[2019]= 16'he60;
assign q[2020]= 16'he85;
assign q[2021]= 16'hebd;
assign q[2022]= 16'hf0c;
assign q[2023]= 16'hf76;
assign q[2024]= 16'hffe;
assign q[2025]= 16'h10a7;
assign q[2026]= 16'h1175;
assign q[2027]= 16'h126b;
assign q[2028]= 16'h1389;
assign q[2029]= 16'h14d2;
assign q[2030]= 16'h1644;
assign q[2031]= 16'h17de;
assign q[2032]= 16'h199f;
assign q[2033]= 16'h1b83;
assign q[2034]= 16'h1d84;
assign q[2035]= 16'h1f9e;
assign q[2036]= 16'h21ca;
assign q[2037]= 16'h2400;
assign q[2038]= 16'h2637;
assign q[2039]= 16'h2866;
assign q[2040]= 16'h2a84;
assign q[2041]= 16'h2c87;
assign q[2042]= 16'h2e64;
assign q[2043]= 16'h3012;
assign q[2044]= 16'h3187;
assign q[2045]= 16'h32bb;
assign q[2046]= 16'h33a3;
assign q[2047]= 16'h343a;
assign q[2048]= 16'h3479;
assign q[2049]= 16'h3459;
assign q[2050]= 16'h33d8;
assign q[2051]= 16'h32f1;
assign q[2052]= 16'h31a2;
assign q[2053]= 16'h2fed;
assign q[2054]= 16'h2dcf;
assign q[2055]= 16'h2b4d;
assign q[2056]= 16'h2867;
assign q[2057]= 16'h2523;
assign q[2058]= 16'h2185;
assign q[2059]= 16'h1d92;
assign q[2060]= 16'h1951;
assign q[2061]= 16'h14c9;
assign q[2062]= 16'h1001;
assign q[2063]= 16'hb04;
assign q[2064]= 16'h5d9;
assign q[2065]= 16'h8b;
assign q[2066]= 16'hfb26;
assign q[2067]= 16'hf5b2;
assign q[2068]= 16'hf03e;
assign q[2069]= 16'head5;
assign q[2070]= 16'he586;
assign q[2071]= 16'he05f;
assign q[2072]= 16'hdb6e;
assign q[2073]= 16'hd6c4;
assign q[2074]= 16'hd26f;
assign q[2075]= 16'hce80;
assign q[2076]= 16'hcb06;
assign q[2077]= 16'hc812;
assign q[2078]= 16'hc5b0;
assign q[2079]= 16'hc3f0;
assign q[2080]= 16'hc2dd;
assign q[2081]= 16'hc281;
assign q[2082]= 16'hc2e4;
assign q[2083]= 16'hc40a;
assign q[2084]= 16'hc5f5;
assign q[2085]= 16'hc8a4;
assign q[2086]= 16'hcc0f;
assign q[2087]= 16'hd02f;
assign q[2088]= 16'hd4f5;
assign q[2089]= 16'hda4f;
assign q[2090]= 16'he028;
assign q[2091]= 16'he667;
assign q[2092]= 16'hecef;
assign q[2093]= 16'hf3a1;
assign q[2094]= 16'hfa5b;
assign q[2095]= 16'hfc;
assign q[2096]= 16'h761;
assign q[2097]= 16'hd66;
assign q[2098]= 16'h12ec;
assign q[2099]= 16'h17d2;
assign q[2100]= 16'h1bfc;
assign q[2101]= 16'h1f53;
assign q[2102]= 16'h21c3;
assign q[2103]= 16'h233e;
assign q[2104]= 16'h23bb;
assign q[2105]= 16'h2337;
assign q[2106]= 16'h21b7;
assign q[2107]= 16'h1f45;
assign q[2108]= 16'h1bf1;
assign q[2109]= 16'h17d1;
assign q[2110]= 16'h12ff;
assign q[2111]= 16'hd9b;
assign q[2112]= 16'h7c6;
assign q[2113]= 16'h1a7;
assign q[2114]= 16'hfb65;
assign q[2115]= 16'hf524;
assign q[2116]= 16'hef0b;
assign q[2117]= 16'he93f;
assign q[2118]= 16'he3e1;
assign q[2119]= 16'hdf0e;
assign q[2120]= 16'hdadf;
assign q[2121]= 16'hd76a;
assign q[2122]= 16'hd4bb;
assign q[2123]= 16'hd2db;
assign q[2124]= 16'hd1cd;
assign q[2125]= 16'hd18e;
assign q[2126]= 16'hd216;
assign q[2127]= 16'hd356;
assign q[2128]= 16'hd53e;
assign q[2129]= 16'hd7b7;
assign q[2130]= 16'hdaab;
assign q[2131]= 16'hddff;
assign q[2132]= 16'he199;
assign q[2133]= 16'he55e;
assign q[2134]= 16'he936;
assign q[2135]= 16'hed08;
assign q[2136]= 16'hf0c0;
assign q[2137]= 16'hf44b;
assign q[2138]= 16'hf79a;
assign q[2139]= 16'hfaa2;
assign q[2140]= 16'hfd5d;
assign q[2141]= 16'hffc6;
assign q[2142]= 16'h1dc;
assign q[2143]= 16'h3a4;
assign q[2144]= 16'h523;
assign q[2145]= 16'h661;
assign q[2146]= 16'h768;
assign q[2147]= 16'h841;
assign q[2148]= 16'h8f7;
assign q[2149]= 16'h995;
assign q[2150]= 16'ha25;
assign q[2151]= 16'haaf;
assign q[2152]= 16'hb3a;
assign q[2153]= 16'hbc9;
assign q[2154]= 16'hc61;
assign q[2155]= 16'hd01;
assign q[2156]= 16'hda9;
assign q[2157]= 16'he54;
assign q[2158]= 16'heff;
assign q[2159]= 16'hfa3;
assign q[2160]= 16'h1039;
assign q[2161]= 16'h10bc;
assign q[2162]= 16'h1123;
assign q[2163]= 16'h116a;
assign q[2164]= 16'h118c;
assign q[2165]= 16'h1184;
assign q[2166]= 16'h1153;
assign q[2167]= 16'h10f7;
assign q[2168]= 16'h1075;
assign q[2169]= 16'hfd0;
assign q[2170]= 16'hf0f;
assign q[2171]= 16'he3b;
assign q[2172]= 16'hd5d;
assign q[2173]= 16'hc82;
assign q[2174]= 16'hbb4;
assign q[2175]= 16'haff;
assign q[2176]= 16'ha71;
assign q[2177]= 16'ha12;
assign q[2178]= 16'h9ee;
assign q[2179]= 16'ha0d;
assign q[2180]= 16'ha74;
assign q[2181]= 16'hb27;
assign q[2182]= 16'hc28;
assign q[2183]= 16'hd75;
assign q[2184]= 16'hf0a;
assign q[2185]= 16'h10e0;
assign q[2186]= 16'h12ee;
assign q[2187]= 16'h1528;
assign q[2188]= 16'h1783;
assign q[2189]= 16'h19ee;
assign q[2190]= 16'h1c5a;
assign q[2191]= 16'h1eb6;
assign q[2192]= 16'h20f4;
assign q[2193]= 16'h2301;
assign q[2194]= 16'h24d1;
assign q[2195]= 16'h2653;
assign q[2196]= 16'h277e;
assign q[2197]= 16'h2845;
assign q[2198]= 16'h28a1;
assign q[2199]= 16'h288d;
assign q[2200]= 16'h2805;
assign q[2201]= 16'h2707;
assign q[2202]= 16'h2597;
assign q[2203]= 16'h23b6;
assign q[2204]= 16'h216d;
assign q[2205]= 16'h1ec2;
assign q[2206]= 16'h1bc0;
assign q[2207]= 16'h1872;
assign q[2208]= 16'h14e5;
assign q[2209]= 16'h1125;
assign q[2210]= 16'hd42;
assign q[2211]= 16'h949;
assign q[2212]= 16'h54a;
assign q[2213]= 16'h153;
assign q[2214]= 16'hfd73;
assign q[2215]= 16'hf9b8;
assign q[2216]= 16'hf62e;
assign q[2217]= 16'hf2e3;
assign q[2218]= 16'hefe2;
assign q[2219]= 16'hed37;
assign q[2220]= 16'heaea;
assign q[2221]= 16'he904;
assign q[2222]= 16'he78c;
assign q[2223]= 16'he688;
assign q[2224]= 16'he5fd;
assign q[2225]= 16'he5ec;
assign q[2226]= 16'he657;
assign q[2227]= 16'he73d;
assign q[2228]= 16'he89c;
assign q[2229]= 16'hea71;
assign q[2230]= 16'hecb4;
assign q[2231]= 16'hef5f;
assign q[2232]= 16'hf268;
assign q[2233]= 16'hf5c3;
assign q[2234]= 16'hf966;
assign q[2235]= 16'hfd41;
assign q[2236]= 16'h144;
assign q[2237]= 16'h562;
assign q[2238]= 16'h988;
assign q[2239]= 16'hda6;
assign q[2240]= 16'h11ab;
assign q[2241]= 16'h1585;
assign q[2242]= 16'h1926;
assign q[2243]= 16'h1c7d;
assign q[2244]= 16'h1f7d;
assign q[2245]= 16'h221b;
assign q[2246]= 16'h244d;
assign q[2247]= 16'h260b;
assign q[2248]= 16'h2752;
assign q[2249]= 16'h281e;
assign q[2250]= 16'h2871;
assign q[2251]= 16'h284e;
assign q[2252]= 16'h27bb;
assign q[2253]= 16'h26c2;
assign q[2254]= 16'h256c;
assign q[2255]= 16'h23c6;
assign q[2256]= 16'h21e0;
assign q[2257]= 16'h1fc9;
assign q[2258]= 16'h1d91;
assign q[2259]= 16'h1b49;
assign q[2260]= 16'h1901;
assign q[2261]= 16'h16c9;
assign q[2262]= 16'h14ae;
assign q[2263]= 16'h12bf;
assign q[2264]= 16'h1104;
assign q[2265]= 16'hf86;
assign q[2266]= 16'he4c;
assign q[2267]= 16'hd57;
assign q[2268]= 16'hca8;
assign q[2269]= 16'hc3c;
assign q[2270]= 16'hc0e;
assign q[2271]= 16'hc16;
assign q[2272]= 16'hc4a;
assign q[2273]= 16'hc9f;
assign q[2274]= 16'hd08;
assign q[2275]= 16'hd77;
assign q[2276]= 16'hddf;
assign q[2277]= 16'he32;
assign q[2278]= 16'he64;
assign q[2279]= 16'he69;
assign q[2280]= 16'he37;
assign q[2281]= 16'hdc6;
assign q[2282]= 16'hd12;
assign q[2283]= 16'hc17;
assign q[2284]= 16'had6;
assign q[2285]= 16'h951;
assign q[2286]= 16'h78e;
assign q[2287]= 16'h594;
assign q[2288]= 16'h36d;
assign q[2289]= 16'h125;
assign q[2290]= 16'hfec9;
assign q[2291]= 16'hfc66;
assign q[2292]= 16'hfa0a;
assign q[2293]= 16'hf7c3;
assign q[2294]= 16'hf59f;
assign q[2295]= 16'hf3a9;
assign q[2296]= 16'hf1ec;
assign q[2297]= 16'hf06f;
assign q[2298]= 16'hef38;
assign q[2299]= 16'hee4b;
assign q[2300]= 16'hedaa;
assign q[2301]= 16'hed51;
assign q[2302]= 16'hed3d;
assign q[2303]= 16'hed69;
assign q[2304]= 16'hedcb;
assign q[2305]= 16'hee5c;
assign q[2306]= 16'hef10;
assign q[2307]= 16'hefdf;
assign q[2308]= 16'hf0bc;
assign q[2309]= 16'hf1a0;
assign q[2310]= 16'hf283;
assign q[2311]= 16'hf35d;
assign q[2312]= 16'hf42c;
assign q[2313]= 16'hf4ed;
assign q[2314]= 16'hf5a0;
assign q[2315]= 16'hf64a;
assign q[2316]= 16'hf6f0;
assign q[2317]= 16'hf799;
assign q[2318]= 16'hf850;
assign q[2319]= 16'hf920;
assign q[2320]= 16'hfa14;
assign q[2321]= 16'hfb39;
assign q[2322]= 16'hfc99;
assign q[2323]= 16'hfe40;
assign q[2324]= 16'h33;
assign q[2325]= 16'h27b;
assign q[2326]= 16'h518;
assign q[2327]= 16'h809;
assign q[2328]= 16'hb49;
assign q[2329]= 16'hecd;
assign q[2330]= 16'h1289;
assign q[2331]= 16'h166a;
assign q[2332]= 16'h1a5a;
assign q[2333]= 16'h1e41;
assign q[2334]= 16'h2205;
assign q[2335]= 16'h2588;
assign q[2336]= 16'h28ad;
assign q[2337]= 16'h2b59;
assign q[2338]= 16'h2d6e;
assign q[2339]= 16'h2ed5;
assign q[2340]= 16'h2f7a;
assign q[2341]= 16'h2f4b;
assign q[2342]= 16'h2e3d;
assign q[2343]= 16'h2c4d;
assign q[2344]= 16'h297b;
assign q[2345]= 16'h25d0;
assign q[2346]= 16'h215b;
assign q[2347]= 16'h1c34;
assign q[2348]= 16'h1675;
assign q[2349]= 16'h1040;
assign q[2350]= 16'h9bd;
assign q[2351]= 16'h314;
assign q[2352]= 16'hfc72;
assign q[2353]= 16'hf603;
assign q[2354]= 16'heff4;
assign q[2355]= 16'hea6f;
assign q[2356]= 16'he59b;
assign q[2357]= 16'he19c;
assign q[2358]= 16'hde8d;
assign q[2359]= 16'hdc85;
assign q[2360]= 16'hdb93;
assign q[2361]= 16'hdbbd;
assign q[2362]= 16'hdd01;
assign q[2363]= 16'hdf57;
assign q[2364]= 16'he2ad;
assign q[2365]= 16'he6ea;
assign q[2366]= 16'hebee;
assign q[2367]= 16'hf196;
assign q[2368]= 16'hf7b8;
assign q[2369]= 16'hfe29;
assign q[2370]= 16'h4bb;
assign q[2371]= 16'hb43;
assign q[2372]= 16'h1194;
assign q[2373]= 16'h1786;
assign q[2374]= 16'h1cf4;
assign q[2375]= 16'h21be;
assign q[2376]= 16'h25cb;
assign q[2377]= 16'h2908;
assign q[2378]= 16'h2b6a;
assign q[2379]= 16'h2ced;
assign q[2380]= 16'h2d92;
assign q[2381]= 16'h2d63;
assign q[2382]= 16'h2c70;
assign q[2383]= 16'h2acf;
assign q[2384]= 16'h2897;
assign q[2385]= 16'h25e7;
assign q[2386]= 16'h22de;
assign q[2387]= 16'h1f9b;
assign q[2388]= 16'h1c3f;
assign q[2389]= 16'h18e8;
assign q[2390]= 16'h15b3;
assign q[2391]= 16'h12b8;
assign q[2392]= 16'h100c;
assign q[2393]= 16'hdc1;
assign q[2394]= 16'hbe1;
assign q[2395]= 16'ha72;
assign q[2396]= 16'h976;
assign q[2397]= 16'h8e9;
assign q[2398]= 16'h8c3;
assign q[2399]= 16'h8f8;
assign q[2400]= 16'h977;
assign q[2401]= 16'ha30;
assign q[2402]= 16'hb0f;
assign q[2403]= 16'hbff;
assign q[2404]= 16'hcec;
assign q[2405]= 16'hdc4;
assign q[2406]= 16'he73;
assign q[2407]= 16'heea;
assign q[2408]= 16'hf1d;
assign q[2409]= 16'hf02;
assign q[2410]= 16'he92;
assign q[2411]= 16'hdca;
assign q[2412]= 16'hcab;
assign q[2413]= 16'hb38;
assign q[2414]= 16'h978;
assign q[2415]= 16'h772;
assign q[2416]= 16'h532;
assign q[2417]= 16'h2c3;
assign q[2418]= 16'h33;
assign q[2419]= 16'hfd8f;
assign q[2420]= 16'hfae3;
assign q[2421]= 16'hf83a;
assign q[2422]= 16'hf5a0;
assign q[2423]= 16'hf31e;
assign q[2424]= 16'hf0ba;
assign q[2425]= 16'hee79;
assign q[2426]= 16'hec5e;
assign q[2427]= 16'hea6a;
assign q[2428]= 16'he89b;
assign q[2429]= 16'he6ee;
assign q[2430]= 16'he55f;
assign q[2431]= 16'he3e6;
assign q[2432]= 16'he27f;
assign q[2433]= 16'he122;
assign q[2434]= 16'hdfc9;
assign q[2435]= 16'hde6e;
assign q[2436]= 16'hdd0b;
assign q[2437]= 16'hdb9e;
assign q[2438]= 16'hda24;
assign q[2439]= 16'hd89e;
assign q[2440]= 16'hd70c;
assign q[2441]= 16'hd575;
assign q[2442]= 16'hd3dd;
assign q[2443]= 16'hd24d;
assign q[2444]= 16'hd0ce;
assign q[2445]= 16'hcf6b;
assign q[2446]= 16'hce32;
assign q[2447]= 16'hcd2d;
assign q[2448]= 16'hcc6b;
assign q[2449]= 16'hcbf8;
assign q[2450]= 16'hcbde;
assign q[2451]= 16'hcc29;
assign q[2452]= 16'hcce0;
assign q[2453]= 16'hce0a;
assign q[2454]= 16'hcfaa;
assign q[2455]= 16'hd1c0;
assign q[2456]= 16'hd44a;
assign q[2457]= 16'hd741;
assign q[2458]= 16'hda9d;
assign q[2459]= 16'hde50;
assign q[2460]= 16'he24b;
assign q[2461]= 16'he67d;
assign q[2462]= 16'head1;
assign q[2463]= 16'hef32;
assign q[2464]= 16'hf388;
assign q[2465]= 16'hf7bd;
assign q[2466]= 16'hfbb9;
assign q[2467]= 16'hff68;
assign q[2468]= 16'h2b3;
assign q[2469]= 16'h58b;
assign q[2470]= 16'h7e1;
assign q[2471]= 16'h9a9;
assign q[2472]= 16'hadc;
assign q[2473]= 16'hb78;
assign q[2474]= 16'hb7f;
assign q[2475]= 16'haf6;
assign q[2476]= 16'h9e9;
assign q[2477]= 16'h867;
assign q[2478]= 16'h682;
assign q[2479]= 16'h44f;
assign q[2480]= 16'h1e8;
assign q[2481]= 16'hff66;
assign q[2482]= 16'hfce3;
assign q[2483]= 16'hfa7a;
assign q[2484]= 16'hf843;
assign q[2485]= 16'hf657;
assign q[2486]= 16'hf4c9;
assign q[2487]= 16'hf3ab;
assign q[2488]= 16'hf308;
assign q[2489]= 16'hf2e8;
assign q[2490]= 16'hf34e;
assign q[2491]= 16'hf437;
assign q[2492]= 16'hf59a;
assign q[2493]= 16'hf76a;
assign q[2494]= 16'hf996;
assign q[2495]= 16'hfc08;
assign q[2496]= 16'hfea8;
assign q[2497]= 16'h15a;
assign q[2498]= 16'h404;
assign q[2499]= 16'h68a;
assign q[2500]= 16'h8d2;
assign q[2501]= 16'hac3;
assign q[2502]= 16'hc47;
assign q[2503]= 16'hd4f;
assign q[2504]= 16'hdcf;
assign q[2505]= 16'hdc0;
assign q[2506]= 16'hd21;
assign q[2507]= 16'hbf7;
assign q[2508]= 16'ha4f;
assign q[2509]= 16'h837;
assign q[2510]= 16'h5c6;
assign q[2511]= 16'h315;
assign q[2512]= 16'h3f;
assign q[2513]= 16'hfd63;
assign q[2514]= 16'hfa9f;
assign q[2515]= 16'hf811;
assign q[2516]= 16'hf5d5;
assign q[2517]= 16'hf404;
assign q[2518]= 16'hf2b2;
assign q[2519]= 16'hf1ef;
assign q[2520]= 16'hf1c5;
assign q[2521]= 16'hf236;
assign q[2522]= 16'hf340;
assign q[2523]= 16'hf4d7;
assign q[2524]= 16'hf6ed;
assign q[2525]= 16'hf969;
assign q[2526]= 16'hfc33;
assign q[2527]= 16'hff2a;
assign q[2528]= 16'h22c;
assign q[2529]= 16'h519;
assign q[2530]= 16'h7cc;
assign q[2531]= 16'ha24;
assign q[2532]= 16'hc03;
assign q[2533]= 16'hd4f;
assign q[2534]= 16'hdf2;
assign q[2535]= 16'hddd;
assign q[2536]= 16'hd09;
assign q[2537]= 16'hb74;
assign q[2538]= 16'h925;
assign q[2539]= 16'h629;
assign q[2540]= 16'h295;
assign q[2541]= 16'hfe85;
assign q[2542]= 16'hfa15;
assign q[2543]= 16'hf56a;
assign q[2544]= 16'hf0a9;
assign q[2545]= 16'hebfb;
assign q[2546]= 16'he785;
assign q[2547]= 16'he36c;
assign q[2548]= 16'hdfd3;
assign q[2549]= 16'hdcd7;
assign q[2550]= 16'hda91;
assign q[2551]= 16'hd912;
assign q[2552]= 16'hd866;
assign q[2553]= 16'hd890;
assign q[2554]= 16'hd98e;
assign q[2555]= 16'hdb55;
assign q[2556]= 16'hddd4;
assign q[2557]= 16'he0f5;
assign q[2558]= 16'he49b;
assign q[2559]= 16'he8a7;
assign q[2560]= 16'hecf7;
assign q[2561]= 16'hf165;
assign q[2562]= 16'hf5ce;
assign q[2563]= 16'hfa0d;
assign q[2564]= 16'hfe02;
assign q[2565]= 16'h18b;
assign q[2566]= 16'h491;
assign q[2567]= 16'h6fb;
assign q[2568]= 16'h8ba;
assign q[2569]= 16'h9c0;
assign q[2570]= 16'ha08;
assign q[2571]= 16'h990;
assign q[2572]= 16'h85d;
assign q[2573]= 16'h678;
assign q[2574]= 16'h3ed;
assign q[2575]= 16'hcd;
assign q[2576]= 16'hfd2d;
assign q[2577]= 16'hf920;
assign q[2578]= 16'hf4bf;
assign q[2579]= 16'hf020;
assign q[2580]= 16'heb5d;
assign q[2581]= 16'he68d;
assign q[2582]= 16'he1c7;
assign q[2583]= 16'hdd20;
assign q[2584]= 16'hd8ae;
assign q[2585]= 16'hd484;
assign q[2586]= 16'hd0b2;
assign q[2587]= 16'hcd47;
assign q[2588]= 16'hca53;
assign q[2589]= 16'hc7e0;
assign q[2590]= 16'hc5fa;
assign q[2591]= 16'hc4a9;
assign q[2592]= 16'hc3f4;
assign q[2593]= 16'hc3e1;
assign q[2594]= 16'hc473;
assign q[2595]= 16'hc5ad;
assign q[2596]= 16'hc78f;
assign q[2597]= 16'hca15;
assign q[2598]= 16'hcd3d;
assign q[2599]= 16'hd0fd;
assign q[2600]= 16'hd54e;
assign q[2601]= 16'hda22;
assign q[2602]= 16'hdf6a;
assign q[2603]= 16'he513;
assign q[2604]= 16'heb0a;
assign q[2605]= 16'hf138;
assign q[2606]= 16'hf782;
assign q[2607]= 16'hfdd0;
assign q[2608]= 16'h404;
assign q[2609]= 16'ha04;
assign q[2610]= 16'hfb5;
assign q[2611]= 16'h14fe;
assign q[2612]= 16'h19c5;
assign q[2613]= 16'h1df6;
assign q[2614]= 16'h2181;
assign q[2615]= 16'h2459;
assign q[2616]= 16'h2674;
assign q[2617]= 16'h27d2;
assign q[2618]= 16'h2873;
assign q[2619]= 16'h2862;
assign q[2620]= 16'h27ab;
assign q[2621]= 16'h2661;
assign q[2622]= 16'h249a;
assign q[2623]= 16'h2272;
assign q[2624]= 16'h2005;
assign q[2625]= 16'h1d72;
assign q[2626]= 16'h1ad9;
assign q[2627]= 16'h1859;
assign q[2628]= 16'h160f;
assign q[2629]= 16'h1416;
assign q[2630]= 16'h1284;
assign q[2631]= 16'h116b;
assign q[2632]= 16'h10d7;
assign q[2633]= 16'h10cf;
assign q[2634]= 16'h1155;
assign q[2635]= 16'h1261;
assign q[2636]= 16'h13ea;
assign q[2637]= 16'h15dd;
assign q[2638]= 16'h1826;
assign q[2639]= 16'h1aaa;
assign q[2640]= 16'h1d4d;
assign q[2641]= 16'h1ff2;
assign q[2642]= 16'h2278;
assign q[2643]= 16'h24c3;
assign q[2644]= 16'h26b6;
assign q[2645]= 16'h2837;
assign q[2646]= 16'h2932;
assign q[2647]= 16'h2996;
assign q[2648]= 16'h2957;
assign q[2649]= 16'h2871;
assign q[2650]= 16'h26e3;
assign q[2651]= 16'h24b5;
assign q[2652]= 16'h21f2;
assign q[2653]= 16'h1eac;
assign q[2654]= 16'h1af9;
assign q[2655]= 16'h16f1;
assign q[2656]= 16'h12b1;
assign q[2657]= 16'he56;
assign q[2658]= 16'h9fe;
assign q[2659]= 16'h5c6;
assign q[2660]= 16'h1cb;
assign q[2661]= 16'hfe27;
assign q[2662]= 16'hfaed;
assign q[2663]= 16'hf831;
assign q[2664]= 16'hf601;
assign q[2665]= 16'hf465;
assign q[2666]= 16'hf362;
assign q[2667]= 16'hf2f7;
assign q[2668]= 16'hf31e;
assign q[2669]= 16'hf3ce;
assign q[2670]= 16'hf4fb;
assign q[2671]= 16'hf694;
assign q[2672]= 16'hf886;
assign q[2673]= 16'hfabd;
assign q[2674]= 16'hfd25;
assign q[2675]= 16'hffa6;
assign q[2676]= 16'h22c;
assign q[2677]= 16'h4a3;
assign q[2678]= 16'h6f8;
assign q[2679]= 16'h918;
assign q[2680]= 16'haf5;
assign q[2681]= 16'hc80;
assign q[2682]= 16'hdb0;
assign q[2683]= 16'he7a;
assign q[2684]= 16'hed9;
assign q[2685]= 16'hec8;
assign q[2686]= 16'he45;
assign q[2687]= 16'hd4f;
assign q[2688]= 16'hbe8;
assign q[2689]= 16'ha13;
assign q[2690]= 16'h7d4;
assign q[2691]= 16'h532;
assign q[2692]= 16'h235;
assign q[2693]= 16'hfee7;
assign q[2694]= 16'hfb50;
assign q[2695]= 16'hf77f;
assign q[2696]= 16'hf381;
assign q[2697]= 16'hef66;
assign q[2698]= 16'heb40;
assign q[2699]= 16'he720;
assign q[2700]= 16'he31b;
assign q[2701]= 16'hdf46;
assign q[2702]= 16'hdbb6;
assign q[2703]= 16'hd881;
assign q[2704]= 16'hd5bc;
assign q[2705]= 16'hd37d;
assign q[2706]= 16'hd1d7;
assign q[2707]= 16'hd0db;
assign q[2708]= 16'hd096;
assign q[2709]= 16'hd116;
assign q[2710]= 16'hd25f;
assign q[2711]= 16'hd475;
assign q[2712]= 16'hd754;
assign q[2713]= 16'hdaf6;
assign q[2714]= 16'hdf4c;
assign q[2715]= 16'he443;
assign q[2716]= 16'he9c4;
assign q[2717]= 16'hefb2;
assign q[2718]= 16'hf5ed;
assign q[2719]= 16'hfc51;
assign q[2720]= 16'h2b7;
assign q[2721]= 16'h8fa;
assign q[2722]= 16'hef1;
assign q[2723]= 16'h1477;
assign q[2724]= 16'h1969;
assign q[2725]= 16'h1da7;
assign q[2726]= 16'h2116;
assign q[2727]= 16'h23a3;
assign q[2728]= 16'h253f;
assign q[2729]= 16'h25e3;
assign q[2730]= 16'h2590;
assign q[2731]= 16'h244f;
assign q[2732]= 16'h2231;
assign q[2733]= 16'h1f4c;
assign q[2734]= 16'h1bbf;
assign q[2735]= 16'h17ae;
assign q[2736]= 16'h133e;
assign q[2737]= 16'he9d;
assign q[2738]= 16'h9f4;
assign q[2739]= 16'h571;
assign q[2740]= 16'h13f;
assign q[2741]= 16'hfd85;
assign q[2742]= 16'hfa65;
assign q[2743]= 16'hf7fe;
assign q[2744]= 16'hf667;
assign q[2745]= 16'hf5ae;
assign q[2746]= 16'hf5dc;
assign q[2747]= 16'hf6ef;
assign q[2748]= 16'hf8df;
assign q[2749]= 16'hfb9a;
assign q[2750]= 16'hff08;
assign q[2751]= 16'h309;
assign q[2752]= 16'h77d;
assign q[2753]= 16'hc39;
assign q[2754]= 16'h1115;
assign q[2755]= 16'h15e5;
assign q[2756]= 16'h1a7e;
assign q[2757]= 16'h1eb8;
assign q[2758]= 16'h226d;
assign q[2759]= 16'h257d;
assign q[2760]= 16'h27cc;
assign q[2761]= 16'h2947;
assign q[2762]= 16'h29e0;
assign q[2763]= 16'h2991;
assign q[2764]= 16'h285b;
assign q[2765]= 16'h2647;
assign q[2766]= 16'h2364;
assign q[2767]= 16'h1fc7;
assign q[2768]= 16'h1b89;
assign q[2769]= 16'h16ca;
assign q[2770]= 16'h11a8;
assign q[2771]= 16'hc47;
assign q[2772]= 16'h6c8;
assign q[2773]= 16'h14c;
assign q[2774]= 16'hfbf3;
assign q[2775]= 16'hf6d6;
assign q[2776]= 16'hf20e;
assign q[2777]= 16'hedad;
assign q[2778]= 16'he9c2;
assign q[2779]= 16'he653;
assign q[2780]= 16'he366;
assign q[2781]= 16'he0f6;
assign q[2782]= 16'hdeff;
assign q[2783]= 16'hdd76;
assign q[2784]= 16'hdc4e;
assign q[2785]= 16'hdb78;
assign q[2786]= 16'hdae2;
assign q[2787]= 16'hda7d;
assign q[2788]= 16'hda39;
assign q[2789]= 16'hda07;
assign q[2790]= 16'hd9dc;
assign q[2791]= 16'hd9af;
assign q[2792]= 16'hd97c;
assign q[2793]= 16'hd941;
assign q[2794]= 16'hd901;
assign q[2795]= 16'hd8c2;
assign q[2796]= 16'hd88f;
assign q[2797]= 16'hd876;
assign q[2798]= 16'hd884;
assign q[2799]= 16'hd8cb;
assign q[2800]= 16'hd95c;
assign q[2801]= 16'hda49;
assign q[2802]= 16'hdba0;
assign q[2803]= 16'hdd70;
assign q[2804]= 16'hdfc2;
assign q[2805]= 16'he29d;
assign q[2806]= 16'he601;
assign q[2807]= 16'he9ec;
assign q[2808]= 16'hee56;
assign q[2809]= 16'hf330;
assign q[2810]= 16'hf867;
assign q[2811]= 16'hfde3;
assign q[2812]= 16'h388;
assign q[2813]= 16'h938;
assign q[2814]= 16'hed2;
assign q[2815]= 16'h1430;
assign q[2816]= 16'h1932;
assign q[2817]= 16'h1db3;
assign q[2818]= 16'h2195;
assign q[2819]= 16'h24ba;
assign q[2820]= 16'h270a;
assign q[2821]= 16'h2871;
assign q[2822]= 16'h28e3;
assign q[2823]= 16'h2859;
assign q[2824]= 16'h26d3;
assign q[2825]= 16'h2458;
assign q[2826]= 16'h20f8;
assign q[2827]= 16'h1cc7;
assign q[2828]= 16'h17e1;
assign q[2829]= 16'h1267;
assign q[2830]= 16'hc7d;
assign q[2831]= 16'h64d;
assign q[2832]= 16'h1;
assign q[2833]= 16'hf9c7;
assign q[2834]= 16'hf3c6;
assign q[2835]= 16'hee2c;
assign q[2836]= 16'he91d;
assign q[2837]= 16'he4bf;
assign q[2838]= 16'he130;
assign q[2839]= 16'hde87;
assign q[2840]= 16'hdcd8;
assign q[2841]= 16'hdc2f;
assign q[2842]= 16'hdc90;
assign q[2843]= 16'hddf9;
assign q[2844]= 16'he061;
assign q[2845]= 16'he3ba;
assign q[2846]= 16'he7ee;
assign q[2847]= 16'hece3;
assign q[2848]= 16'hf27c;
assign q[2849]= 16'hf896;
assign q[2850]= 16'hff0e;
assign q[2851]= 16'h5c0;
assign q[2852]= 16'hc86;
assign q[2853]= 16'h133e;
assign q[2854]= 16'h19c3;
assign q[2855]= 16'h1ff6;
assign q[2856]= 16'h25bc;
assign q[2857]= 16'h2afa;
assign q[2858]= 16'h2f9c;
assign q[2859]= 16'h3392;
assign q[2860]= 16'h36d0;
assign q[2861]= 16'h3950;
assign q[2862]= 16'h3b0e;
assign q[2863]= 16'h3c0d;
assign q[2864]= 16'h3c51;
assign q[2865]= 16'h3be4;
assign q[2866]= 16'h3ad1;
assign q[2867]= 16'h3926;
assign q[2868]= 16'h36f2;
assign q[2869]= 16'h3447;
assign q[2870]= 16'h3136;
assign q[2871]= 16'h2dd1;
assign q[2872]= 16'h2a2a;
assign q[2873]= 16'h2653;
assign q[2874]= 16'h225c;
assign q[2875]= 16'h1e54;
assign q[2876]= 16'h1a4b;
assign q[2877]= 16'h164c;
assign q[2878]= 16'h1265;
assign q[2879]= 16'he9f;
assign q[2880]= 16'hb04;
assign q[2881]= 16'h79d;
assign q[2882]= 16'h470;
assign q[2883]= 16'h184;
assign q[2884]= 16'hfee0;
assign q[2885]= 16'hfc86;
assign q[2886]= 16'hfa7c;
assign q[2887]= 16'hf8c4;
assign q[2888]= 16'hf761;
assign q[2889]= 16'hf657;
assign q[2890]= 16'hf5a6;
assign q[2891]= 16'hf54f;
assign q[2892]= 16'hf553;
assign q[2893]= 16'hf5b1;
assign q[2894]= 16'hf668;
assign q[2895]= 16'hf775;
assign q[2896]= 16'hf8d4;
assign q[2897]= 16'hfa82;
assign q[2898]= 16'hfc78;
assign q[2899]= 16'hfeb2;
assign q[2900]= 16'h125;
assign q[2901]= 16'h3cb;
assign q[2902]= 16'h69b;
assign q[2903]= 16'h98b;
assign q[2904]= 16'hc8f;
assign q[2905]= 16'hf9e;
assign q[2906]= 16'h12ab;
assign q[2907]= 16'h15ad;
assign q[2908]= 16'h1899;
assign q[2909]= 16'h1b63;
assign q[2910]= 16'h1e02;
assign q[2911]= 16'h206e;
assign q[2912]= 16'h229f;
assign q[2913]= 16'h248d;
assign q[2914]= 16'h2634;
assign q[2915]= 16'h278e;
assign q[2916]= 16'h2898;
assign q[2917]= 16'h2952;
assign q[2918]= 16'h29bb;
assign q[2919]= 16'h29d4;
assign q[2920]= 16'h29a0;
assign q[2921]= 16'h2922;
assign q[2922]= 16'h285e;
assign q[2923]= 16'h275b;
assign q[2924]= 16'h261e;
assign q[2925]= 16'h24b0;
assign q[2926]= 16'h2317;
assign q[2927]= 16'h215b;
assign q[2928]= 16'h1f86;
assign q[2929]= 16'h1d9f;
assign q[2930]= 16'h1baf;
assign q[2931]= 16'h19bd;
assign q[2932]= 16'h17d3;
assign q[2933]= 16'h15f6;
assign q[2934]= 16'h142f;
assign q[2935]= 16'h1283;
assign q[2936]= 16'h10f7;
assign q[2937]= 16'hf92;
assign q[2938]= 16'he56;
assign q[2939]= 16'hd47;
assign q[2940]= 16'hc68;
assign q[2941]= 16'hbb9;
assign q[2942]= 16'hb3c;
assign q[2943]= 16'haf0;
assign q[2944]= 16'had5;
assign q[2945]= 16'haea;
assign q[2946]= 16'hb2c;
assign q[2947]= 16'hb99;
assign q[2948]= 16'hc2e;
assign q[2949]= 16'hce9;
assign q[2950]= 16'hdc7;
assign q[2951]= 16'hec4;
assign q[2952]= 16'hfde;
assign q[2953]= 16'h1111;
assign q[2954]= 16'h125c;
assign q[2955]= 16'h13bb;
assign q[2956]= 16'h152c;
assign q[2957]= 16'h16ae;
assign q[2958]= 16'h183f;
assign q[2959]= 16'h19dd;
assign q[2960]= 16'h1b88;
assign q[2961]= 16'h1d3d;
assign q[2962]= 16'h1efb;
assign q[2963]= 16'h20c1;
assign q[2964]= 16'h228d;
assign q[2965]= 16'h245b;
assign q[2966]= 16'h2628;
assign q[2967]= 16'h27f1;
assign q[2968]= 16'h29b2;
assign q[2969]= 16'h2b63;
assign q[2970]= 16'h2d00;
assign q[2971]= 16'h2e82;
assign q[2972]= 16'h2fe0;
assign q[2973]= 16'h3113;
assign q[2974]= 16'h3213;
assign q[2975]= 16'h32d7;
assign q[2976]= 16'h3356;
assign q[2977]= 16'h338a;
assign q[2978]= 16'h336a;
assign q[2979]= 16'h32f0;
assign q[2980]= 16'h3219;
assign q[2981]= 16'h30e0;
assign q[2982]= 16'h2f44;
assign q[2983]= 16'h2d46;
assign q[2984]= 16'h2ae8;
assign q[2985]= 16'h2830;
assign q[2986]= 16'h2524;
assign q[2987]= 16'h21ce;
assign q[2988]= 16'h1e3a;
assign q[2989]= 16'h1a73;
assign q[2990]= 16'h168a;
assign q[2991]= 16'h128f;
assign q[2992]= 16'he91;
assign q[2993]= 16'haa3;
assign q[2994]= 16'h6d6;
assign q[2995]= 16'h33a;
assign q[2996]= 16'hffe2;
assign q[2997]= 16'hfcd9;
assign q[2998]= 16'hfa2d;
assign q[2999]= 16'hf7ea;
assign q[3000]= 16'hf618;
assign q[3001]= 16'hf4be;
assign q[3002]= 16'hf3df;
assign q[3003]= 16'hf37c;
assign q[3004]= 16'hf393;
assign q[3005]= 16'hf420;
assign q[3006]= 16'hf51e;
assign q[3007]= 16'hf682;
assign q[3008]= 16'hf844;
assign q[3009]= 16'hfa57;
assign q[3010]= 16'hfcaf;
assign q[3011]= 16'hff3f;
assign q[3012]= 16'h1f8;
assign q[3013]= 16'h4d0;
assign q[3014]= 16'h7b8;
assign q[3015]= 16'haa5;
assign q[3016]= 16'hd8b;
assign q[3017]= 16'h1063;
assign q[3018]= 16'h1322;
assign q[3019]= 16'h15c3;
assign q[3020]= 16'h1841;
assign q[3021]= 16'h1a98;
assign q[3022]= 16'h1cc6;
assign q[3023]= 16'h1ec9;
assign q[3024]= 16'h20a3;
assign q[3025]= 16'h2252;
assign q[3026]= 16'h23da;
assign q[3027]= 16'h253d;
assign q[3028]= 16'h267b;
assign q[3029]= 16'h2799;
assign q[3030]= 16'h2899;
assign q[3031]= 16'h297c;
assign q[3032]= 16'h2a45;
assign q[3033]= 16'h2af5;
assign q[3034]= 16'h2b8f;
assign q[3035]= 16'h2c12;
assign q[3036]= 16'h2c80;
assign q[3037]= 16'h2cd9;
assign q[3038]= 16'h2d1e;
assign q[3039]= 16'h2d4e;
assign q[3040]= 16'h2d6a;
assign q[3041]= 16'h2d71;
assign q[3042]= 16'h2d64;
assign q[3043]= 16'h2d43;
assign q[3044]= 16'h2d0c;
assign q[3045]= 16'h2cc2;
assign q[3046]= 16'h2c62;
assign q[3047]= 16'h2bec;
assign q[3048]= 16'h2b61;
assign q[3049]= 16'h2abe;
assign q[3050]= 16'h2a02;
assign q[3051]= 16'h292c;
assign q[3052]= 16'h283a;
assign q[3053]= 16'h2728;
assign q[3054]= 16'h25f3;
assign q[3055]= 16'h2498;
assign q[3056]= 16'h2312;
assign q[3057]= 16'h215e;
assign q[3058]= 16'h1f77;
assign q[3059]= 16'h1d5b;
assign q[3060]= 16'h1b05;
assign q[3061]= 16'h1873;
assign q[3062]= 16'h15a3;
assign q[3063]= 16'h1297;
assign q[3064]= 16'hf4e;
assign q[3065]= 16'hbcb;
assign q[3066]= 16'h815;
assign q[3067]= 16'h430;
assign q[3068]= 16'h27;
assign q[3069]= 16'hfc04;
assign q[3070]= 16'hf7d3;
assign q[3071]= 16'hf3a1;
assign q[3072]= 16'hef7e;
assign q[3073]= 16'heb79;
assign q[3074]= 16'he7a3;
assign q[3075]= 16'he40b;
assign q[3076]= 16'he0c2;
assign q[3077]= 16'hddd6;
assign q[3078]= 16'hdb53;
assign q[3079]= 16'hd944;
assign q[3080]= 16'hd7b1;
assign q[3081]= 16'hd6a1;
assign q[3082]= 16'hd614;
assign q[3083]= 16'hd60c;
assign q[3084]= 16'hd683;
assign q[3085]= 16'hd773;
assign q[3086]= 16'hd8d2;
assign q[3087]= 16'hda94;
assign q[3088]= 16'hdca9;
assign q[3089]= 16'hdf02;
assign q[3090]= 16'he18e;
assign q[3091]= 16'he43a;
assign q[3092]= 16'he6f7;
assign q[3093]= 16'he9b2;
assign q[3094]= 16'hec5e;
assign q[3095]= 16'heeee;
assign q[3096]= 16'hf157;
assign q[3097]= 16'hf393;
assign q[3098]= 16'hf59d;
assign q[3099]= 16'hf774;
assign q[3100]= 16'hf91a;
assign q[3101]= 16'hfa96;
assign q[3102]= 16'hfbef;
assign q[3103]= 16'hfd2f;
assign q[3104]= 16'hfe63;
assign q[3105]= 16'hff97;
assign q[3106]= 16'hd9;
assign q[3107]= 16'h237;
assign q[3108]= 16'h3bc;
assign q[3109]= 16'h572;
assign q[3110]= 16'h761;
assign q[3111]= 16'h98e;
assign q[3112]= 16'hbf8;
assign q[3113]= 16'he9f;
assign q[3114]= 16'h117b;
assign q[3115]= 16'h1483;
assign q[3116]= 16'h17a8;
assign q[3117]= 16'h1ada;
assign q[3118]= 16'h1e05;
assign q[3119]= 16'h2113;
assign q[3120]= 16'h23ee;
assign q[3121]= 16'h267f;
assign q[3122]= 16'h28b0;
assign q[3123]= 16'h2a6b;
assign q[3124]= 16'h2b9e;
assign q[3125]= 16'h2c3b;
assign q[3126]= 16'h2c35;
assign q[3127]= 16'h2b87;
assign q[3128]= 16'h2a2e;
assign q[3129]= 16'h282f;
assign q[3130]= 16'h2593;
assign q[3131]= 16'h2268;
assign q[3132]= 16'h1ec2;
assign q[3133]= 16'h1ab7;
assign q[3134]= 16'h1665;
assign q[3135]= 16'h11e8;
assign q[3136]= 16'hd62;
assign q[3137]= 16'h8f3;
assign q[3138]= 16'h4bd;
assign q[3139]= 16'hde;
assign q[3140]= 16'hfd77;
assign q[3141]= 16'hfa9d;
assign q[3142]= 16'hf869;
assign q[3143]= 16'hf6eb;
assign q[3144]= 16'hf62e;
assign q[3145]= 16'hf638;
assign q[3146]= 16'hf708;
assign q[3147]= 16'hf897;
assign q[3148]= 16'hfada;
assign q[3149]= 16'hfdbe;
assign q[3150]= 16'h12c;
assign q[3151]= 16'h50b;
assign q[3152]= 16'h93e;
assign q[3153]= 16'hda4;
assign q[3154]= 16'h121d;
assign q[3155]= 16'h168a;
assign q[3156]= 16'h1ac9;
assign q[3157]= 16'h1ebf;
assign q[3158]= 16'h2252;
assign q[3159]= 16'h256a;
assign q[3160]= 16'h27f6;
assign q[3161]= 16'h29e8;
assign q[3162]= 16'h2b38;
assign q[3163]= 16'h2be3;
assign q[3164]= 16'h2beb;
assign q[3165]= 16'h2b55;
assign q[3166]= 16'h2a2e;
assign q[3167]= 16'h2884;
assign q[3168]= 16'h2667;
assign q[3169]= 16'h23ec;
assign q[3170]= 16'h2127;
assign q[3171]= 16'h1e2f;
assign q[3172]= 16'h1b18;
assign q[3173]= 16'h17f8;
assign q[3174]= 16'h14df;
assign q[3175]= 16'h11de;
assign q[3176]= 16'hf03;
assign q[3177]= 16'hc57;
assign q[3178]= 16'h9e1;
assign q[3179]= 16'h7a3;
assign q[3180]= 16'h59e;
assign q[3181]= 16'h3cf;
assign q[3182]= 16'h22e;
assign q[3183]= 16'hb4;
assign q[3184]= 16'hff57;
assign q[3185]= 16'hfe0a;
assign q[3186]= 16'hfcc2;
assign q[3187]= 16'hfb73;
assign q[3188]= 16'hfa12;
assign q[3189]= 16'hf896;
assign q[3190]= 16'hf6f6;
assign q[3191]= 16'hf52d;
assign q[3192]= 16'hf338;
assign q[3193]= 16'hf118;
assign q[3194]= 16'heece;
assign q[3195]= 16'hec61;
assign q[3196]= 16'he9d8;
assign q[3197]= 16'he73f;
assign q[3198]= 16'he4a3;
assign q[3199]= 16'he211;
assign q[3200]= 16'hdf9a;
assign q[3201]= 16'hdd4e;
assign q[3202]= 16'hdb3d;
assign q[3203]= 16'hd977;
assign q[3204]= 16'hd80a;
assign q[3205]= 16'hd703;
assign q[3206]= 16'hd66e;
assign q[3207]= 16'hd652;
assign q[3208]= 16'hd6b5;
assign q[3209]= 16'hd79a;
assign q[3210]= 16'hd901;
assign q[3211]= 16'hdae7;
assign q[3212]= 16'hdd45;
assign q[3213]= 16'he014;
assign q[3214]= 16'he348;
assign q[3215]= 16'he6d3;
assign q[3216]= 16'heaa9;
assign q[3217]= 16'heeb8;
assign q[3218]= 16'hf2f1;
assign q[3219]= 16'hf743;
assign q[3220]= 16'hfb9e;
assign q[3221]= 16'hfff2;
assign q[3222]= 16'h430;
assign q[3223]= 16'h84d;
assign q[3224]= 16'hc3c;
assign q[3225]= 16'hff5;
assign q[3226]= 16'h136f;
assign q[3227]= 16'h16a5;
assign q[3228]= 16'h1994;
assign q[3229]= 16'h1c3a;
assign q[3230]= 16'h1e96;
assign q[3231]= 16'h20ab;
assign q[3232]= 16'h227a;
assign q[3233]= 16'h2406;
assign q[3234]= 16'h2555;
assign q[3235]= 16'h2668;
assign q[3236]= 16'h2746;
assign q[3237]= 16'h27f0;
assign q[3238]= 16'h286b;
assign q[3239]= 16'h28b9;
assign q[3240]= 16'h28db;
assign q[3241]= 16'h28d3;
assign q[3242]= 16'h289e;
assign q[3243]= 16'h283e;
assign q[3244]= 16'h27af;
assign q[3245]= 16'h26ef;
assign q[3246]= 16'h25fc;
assign q[3247]= 16'h24d2;
assign q[3248]= 16'h236e;
assign q[3249]= 16'h21cd;
assign q[3250]= 16'h1fee;
assign q[3251]= 16'h1dcf;
assign q[3252]= 16'h1b6f;
assign q[3253]= 16'h18cf;
assign q[3254]= 16'h15f1;
assign q[3255]= 16'h12d7;
assign q[3256]= 16'hf87;
assign q[3257]= 16'hc06;
assign q[3258]= 16'h85b;
assign q[3259]= 16'h48e;
assign q[3260]= 16'ha7;
assign q[3261]= 16'hfcb2;
assign q[3262]= 16'hf8b6;
assign q[3263]= 16'hf4bf;
assign q[3264]= 16'hf0d6;
assign q[3265]= 16'hed05;
assign q[3266]= 16'he956;
assign q[3267]= 16'he5d1;
assign q[3268]= 16'he27e;
assign q[3269]= 16'hdf63;
assign q[3270]= 16'hdc86;
assign q[3271]= 16'hd9eb;
assign q[3272]= 16'hd795;
assign q[3273]= 16'hd587;
assign q[3274]= 16'hd3c0;
assign q[3275]= 16'hd240;
assign q[3276]= 16'hd108;
assign q[3277]= 16'hd014;
assign q[3278]= 16'hcf62;
assign q[3279]= 16'hceef;
assign q[3280]= 16'hceb9;
assign q[3281]= 16'hcebc;
assign q[3282]= 16'hcef4;
assign q[3283]= 16'hcf5e;
assign q[3284]= 16'hcff8;
assign q[3285]= 16'hd0bd;
assign q[3286]= 16'hd1ab;
assign q[3287]= 16'hd2bf;
assign q[3288]= 16'hd3f6;
assign q[3289]= 16'hd54d;
assign q[3290]= 16'hd6c3;
assign q[3291]= 16'hd854;
assign q[3292]= 16'hd9fd;
assign q[3293]= 16'hdbbc;
assign q[3294]= 16'hdd8d;
assign q[3295]= 16'hdf6e;
assign q[3296]= 16'he15b;
assign q[3297]= 16'he350;
assign q[3298]= 16'he54b;
assign q[3299]= 16'he748;
assign q[3300]= 16'he943;
assign q[3301]= 16'heb3a;
assign q[3302]= 16'hed2b;
assign q[3303]= 16'hef13;
assign q[3304]= 16'hf0f0;
assign q[3305]= 16'hf2c3;
assign q[3306]= 16'hf48a;
assign q[3307]= 16'hf645;
assign q[3308]= 16'hf7f7;
assign q[3309]= 16'hf9a1;
assign q[3310]= 16'hfb45;
assign q[3311]= 16'hfce5;
assign q[3312]= 16'hfe83;
assign q[3313]= 16'h22;
assign q[3314]= 16'h1c5;
assign q[3315]= 16'h36e;
assign q[3316]= 16'h51c;
assign q[3317]= 16'h6d0;
assign q[3318]= 16'h88a;
assign q[3319]= 16'ha45;
assign q[3320]= 16'hbff;
assign q[3321]= 16'hdb2;
assign q[3322]= 16'hf58;
assign q[3323]= 16'h10e9;
assign q[3324]= 16'h125c;
assign q[3325]= 16'h13a8;
assign q[3326]= 16'h14c1;
assign q[3327]= 16'h159f;
assign q[3328]= 16'h1635;
assign q[3329]= 16'h167b;
assign q[3330]= 16'h1668;
assign q[3331]= 16'h15f5;
assign q[3332]= 16'h151b;
assign q[3333]= 16'h13d6;
assign q[3334]= 16'h1227;
assign q[3335]= 16'h100d;
assign q[3336]= 16'hd8d;
assign q[3337]= 16'haae;
assign q[3338]= 16'h778;
assign q[3339]= 16'h3f6;
assign q[3340]= 16'h38;
assign q[3341]= 16'hfc4d;
assign q[3342]= 16'hf844;
assign q[3343]= 16'hf432;
assign q[3344]= 16'hf027;
assign q[3345]= 16'hec37;
assign q[3346]= 16'he874;
assign q[3347]= 16'he4f0;
assign q[3348]= 16'he1b9;
assign q[3349]= 16'hdede;
assign q[3350]= 16'hdc69;
assign q[3351]= 16'hda64;
assign q[3352]= 16'hd8d6;
assign q[3353]= 16'hd7c0;
assign q[3354]= 16'hd724;
assign q[3355]= 16'hd700;
assign q[3356]= 16'hd74e;
assign q[3357]= 16'hd808;
assign q[3358]= 16'hd923;
assign q[3359]= 16'hda96;
assign q[3360]= 16'hdc53;
assign q[3361]= 16'hde4d;
assign q[3362]= 16'he076;
assign q[3363]= 16'he2c0;
assign q[3364]= 16'he51c;
assign q[3365]= 16'he77d;
assign q[3366]= 16'he9d6;
assign q[3367]= 16'hec1b;
assign q[3368]= 16'hee42;
assign q[3369]= 16'hf040;
assign q[3370]= 16'hf20d;
assign q[3371]= 16'hf3a3;
assign q[3372]= 16'hf4fc;
assign q[3373]= 16'hf615;
assign q[3374]= 16'hf6eb;
assign q[3375]= 16'hf77c;
assign q[3376]= 16'hf7ca;
assign q[3377]= 16'hf7d5;
assign q[3378]= 16'hf79f;
assign q[3379]= 16'hf72d;
assign q[3380]= 16'hf684;
assign q[3381]= 16'hf5a8;
assign q[3382]= 16'hf4a1;
assign q[3383]= 16'hf377;
assign q[3384]= 16'hf233;
assign q[3385]= 16'hf0de;
assign q[3386]= 16'hef83;
assign q[3387]= 16'hee2d;
assign q[3388]= 16'hece9;
assign q[3389]= 16'hebc2;
assign q[3390]= 16'heac5;
assign q[3391]= 16'he9fd;
assign q[3392]= 16'he978;
assign q[3393]= 16'he93f;
assign q[3394]= 16'he95e;
assign q[3395]= 16'he9db;
assign q[3396]= 16'heabf;
assign q[3397]= 16'hec0e;
assign q[3398]= 16'hedc9;
assign q[3399]= 16'heff0;
assign q[3400]= 16'hf281;
assign q[3401]= 16'hf575;
assign q[3402]= 16'hf8c2;
assign q[3403]= 16'hfc5f;
assign q[3404]= 16'h3a;
assign q[3405]= 16'h445;
assign q[3406]= 16'h86e;
assign q[3407]= 16'hca1;
assign q[3408]= 16'h10c8;
assign q[3409]= 16'h14cf;
assign q[3410]= 16'h18a2;
assign q[3411]= 16'h1c2d;
assign q[3412]= 16'h1f5e;
assign q[3413]= 16'h2227;
assign q[3414]= 16'h247a;
assign q[3415]= 16'h264d;
assign q[3416]= 16'h279b;
assign q[3417]= 16'h2861;
assign q[3418]= 16'h28a1;
assign q[3419]= 16'h285f;
assign q[3420]= 16'h27a4;
assign q[3421]= 16'h267d;
assign q[3422]= 16'h24f8;
assign q[3423]= 16'h2326;
assign q[3424]= 16'h211c;
assign q[3425]= 16'h1eec;
assign q[3426]= 16'h1cac;
assign q[3427]= 16'h1a70;
assign q[3428]= 16'h184d;
assign q[3429]= 16'h1655;
assign q[3430]= 16'h1499;
assign q[3431]= 16'h1328;
assign q[3432]= 16'h120c;
assign q[3433]= 16'h114f;
assign q[3434]= 16'h10f6;
assign q[3435]= 16'h1104;
assign q[3436]= 16'h1177;
assign q[3437]= 16'h124e;
assign q[3438]= 16'h1381;
assign q[3439]= 16'h1509;
assign q[3440]= 16'h16db;
assign q[3441]= 16'h18eb;
assign q[3442]= 16'h1b2d;
assign q[3443]= 16'h1d94;
assign q[3444]= 16'h2011;
assign q[3445]= 16'h2298;
assign q[3446]= 16'h251b;
assign q[3447]= 16'h278d;
assign q[3448]= 16'h29e3;
assign q[3449]= 16'h2c13;
assign q[3450]= 16'h2e13;
assign q[3451]= 16'h2fdb;
assign q[3452]= 16'h3163;
assign q[3453]= 16'h32a5;
assign q[3454]= 16'h339c;
assign q[3455]= 16'h3444;
assign q[3456]= 16'h3499;
assign q[3457]= 16'h3499;
assign q[3458]= 16'h3442;
assign q[3459]= 16'h3393;
assign q[3460]= 16'h328b;
assign q[3461]= 16'h312b;
assign q[3462]= 16'h2f75;
assign q[3463]= 16'h2d6a;
assign q[3464]= 16'h2b0f;
assign q[3465]= 16'h2867;
assign q[3466]= 16'h2577;
assign q[3467]= 16'h2248;
assign q[3468]= 16'h1edf;
assign q[3469]= 16'h1b46;
assign q[3470]= 16'h1788;
assign q[3471]= 16'h13ad;
assign q[3472]= 16'hfc3;
assign q[3473]= 16'hbd4;
assign q[3474]= 16'h7eb;
assign q[3475]= 16'h415;
assign q[3476]= 16'h5c;
assign q[3477]= 16'hfcca;
assign q[3478]= 16'hf966;
assign q[3479]= 16'hf638;
assign q[3480]= 16'hf343;
assign q[3481]= 16'hf08b;
assign q[3482]= 16'hee11;
assign q[3483]= 16'hebd1;
assign q[3484]= 16'he9c9;
assign q[3485]= 16'he7f1;
assign q[3486]= 16'he644;
assign q[3487]= 16'he4b7;
assign q[3488]= 16'he341;
assign q[3489]= 16'he1d7;
assign q[3490]= 16'he070;
assign q[3491]= 16'hdf03;
assign q[3492]= 16'hdd88;
assign q[3493]= 16'hdbf9;
assign q[3494]= 16'hda52;
assign q[3495]= 16'hd893;
assign q[3496]= 16'hd6be;
assign q[3497]= 16'hd4d7;
assign q[3498]= 16'hd2e7;
assign q[3499]= 16'hd0fa;
assign q[3500]= 16'hcf1e;
assign q[3501]= 16'hcd61;
assign q[3502]= 16'hcbd7;
assign q[3503]= 16'hca93;
assign q[3504]= 16'hc9a6;
assign q[3505]= 16'hc926;
assign q[3506]= 16'hc922;
assign q[3507]= 16'hc9ab;
assign q[3508]= 16'hcacd;
assign q[3509]= 16'hcc91;
assign q[3510]= 16'hcefd;
assign q[3511]= 16'hd211;
assign q[3512]= 16'hd5c9;
assign q[3513]= 16'hda1d;
assign q[3514]= 16'hdefe;
assign q[3515]= 16'he45a;
assign q[3516]= 16'hea1a;
assign q[3517]= 16'hf025;
assign q[3518]= 16'hf65b;
assign q[3519]= 16'hfc9e;
assign q[3520]= 16'h2cc;
assign q[3521]= 16'h8c5;
assign q[3522]= 16'he66;
assign q[3523]= 16'h1390;
assign q[3524]= 16'h1826;
assign q[3525]= 16'h1c0c;
assign q[3526]= 16'h1f2d;
assign q[3527]= 16'h2176;
assign q[3528]= 16'h22d9;
assign q[3529]= 16'h234e;
assign q[3530]= 16'h22d2;
assign q[3531]= 16'h2168;
assign q[3532]= 16'h1f16;
assign q[3533]= 16'h1bea;
assign q[3534]= 16'h17f2;
assign q[3535]= 16'h1345;
assign q[3536]= 16'hdfb;
assign q[3537]= 16'h82e;
assign q[3538]= 16'h1fb;
assign q[3539]= 16'hfb82;
assign q[3540]= 16'hf4e0;
assign q[3541]= 16'hee35;
assign q[3542]= 16'he7a0;
assign q[3543]= 16'he13f;
assign q[3544]= 16'hdb2f;
assign q[3545]= 16'hd589;
assign q[3546]= 16'hd065;
assign q[3547]= 16'hcbd9;
assign q[3548]= 16'hc7f7;
assign q[3549]= 16'hc4cd;
assign q[3550]= 16'hc269;
assign q[3551]= 16'hc0d3;
assign q[3552]= 16'hc00f;
assign q[3553]= 16'hc020;
assign q[3554]= 16'hc105;
assign q[3555]= 16'hc2b8;
assign q[3556]= 16'hc533;
assign q[3557]= 16'hc869;
assign q[3558]= 16'hcc4e;
assign q[3559]= 16'hd0d1;
assign q[3560]= 16'hd5de;
assign q[3561]= 16'hdb61;
assign q[3562]= 16'he143;
assign q[3563]= 16'he76a;
assign q[3564]= 16'hedbd;
assign q[3565]= 16'hf421;
assign q[3566]= 16'hfa7b;
assign q[3567]= 16'hb0;
assign q[3568]= 16'h6a6;
assign q[3569]= 16'hc44;
assign q[3570]= 16'h1172;
assign q[3571]= 16'h161c;
assign q[3572]= 16'h1a2e;
assign q[3573]= 16'h1d9a;
assign q[3574]= 16'h2052;
assign q[3575]= 16'h2250;
assign q[3576]= 16'h238d;
assign q[3577]= 16'h240b;
assign q[3578]= 16'h23cc;
assign q[3579]= 16'h22d9;
assign q[3580]= 16'h213d;
assign q[3581]= 16'h1f06;
assign q[3582]= 16'h1c48;
assign q[3583]= 16'h1916;
assign q[3584]= 16'h1588;
assign q[3585]= 16'h11b7;
assign q[3586]= 16'hdbb;
assign q[3587]= 16'h9b0;
assign q[3588]= 16'h5ae;
assign q[3589]= 16'h1cf;
assign q[3590]= 16'hfe2b;
assign q[3591]= 16'hfad5;
assign q[3592]= 16'hf7e1;
assign q[3593]= 16'hf561;
assign q[3594]= 16'hf361;
assign q[3595]= 16'hf1ec;
assign q[3596]= 16'hf108;
assign q[3597]= 16'hf0b9;
assign q[3598]= 16'hf0ff;
assign q[3599]= 16'hf1d8;
assign q[3600]= 16'hf33e;
assign q[3601]= 16'hf527;
assign q[3602]= 16'hf789;
assign q[3603]= 16'hfa57;
assign q[3604]= 16'hfd81;
assign q[3605]= 16'hf7;
assign q[3606]= 16'h4a9;
assign q[3607]= 16'h884;
assign q[3608]= 16'hc75;
assign q[3609]= 16'h106b;
assign q[3610]= 16'h1453;
assign q[3611]= 16'h181c;
assign q[3612]= 16'h1bb5;
assign q[3613]= 16'h1f0f;
assign q[3614]= 16'h221d;
assign q[3615]= 16'h24d1;
assign q[3616]= 16'h2723;
assign q[3617]= 16'h2909;
assign q[3618]= 16'h2a7e;
assign q[3619]= 16'h2b7f;
assign q[3620]= 16'h2c09;
assign q[3621]= 16'h2c1f;
assign q[3622]= 16'h2bc4;
assign q[3623]= 16'h2afe;
assign q[3624]= 16'h29d6;
assign q[3625]= 16'h2858;
assign q[3626]= 16'h268f;
assign q[3627]= 16'h248b;
assign q[3628]= 16'h225c;
assign q[3629]= 16'h2012;
assign q[3630]= 16'h1dc1;
assign q[3631]= 16'h1b79;
assign q[3632]= 16'h194d;
assign q[3633]= 16'h174d;
assign q[3634]= 16'h1589;
assign q[3635]= 16'h140f;
assign q[3636]= 16'h12eb;
assign q[3637]= 16'h1226;
assign q[3638]= 16'h11c5;
assign q[3639]= 16'h11cc;
assign q[3640]= 16'h1239;
assign q[3641]= 16'h130a;
assign q[3642]= 16'h1437;
assign q[3643]= 16'h15b5;
assign q[3644]= 16'h1777;
assign q[3645]= 16'h196d;
assign q[3646]= 16'h1b84;
assign q[3647]= 16'h1da9;
assign q[3648]= 16'h1fc6;
assign q[3649]= 16'h21c5;
assign q[3650]= 16'h2392;
assign q[3651]= 16'h2518;
assign q[3652]= 16'h2642;
assign q[3653]= 16'h26ff;
assign q[3654]= 16'h2741;
assign q[3655]= 16'h26f9;
assign q[3656]= 16'h2620;
assign q[3657]= 16'h24ae;
assign q[3658]= 16'h22a1;
assign q[3659]= 16'h1ff9;
assign q[3660]= 16'h1cbb;
assign q[3661]= 16'h18ed;
assign q[3662]= 16'h149a;
assign q[3663]= 16'hfcf;
assign q[3664]= 16'ha9b;
assign q[3665]= 16'h510;
assign q[3666]= 16'hff42;
assign q[3667]= 16'hf943;
assign q[3668]= 16'hf32b;
assign q[3669]= 16'hed0e;
assign q[3670]= 16'he704;
assign q[3671]= 16'he122;
assign q[3672]= 16'hdb7f;
assign q[3673]= 16'hd630;
assign q[3674]= 16'hd149;
assign q[3675]= 16'hccde;
assign q[3676]= 16'hc901;
assign q[3677]= 16'hc5c2;
assign q[3678]= 16'hc331;
assign q[3679]= 16'hc159;
assign q[3680]= 16'hc046;
assign q[3681]= 16'hc001;
assign q[3682]= 16'hc08d;
assign q[3683]= 16'hc1ee;
assign q[3684]= 16'hc423;
assign q[3685]= 16'hc728;
assign q[3686]= 16'hcaf3;
assign q[3687]= 16'hcf7a;
assign q[3688]= 16'hd4ab;
assign q[3689]= 16'hda74;
assign q[3690]= 16'he0bb;
assign q[3691]= 16'he766;
assign q[3692]= 16'hee56;
assign q[3693]= 16'hf567;
assign q[3694]= 16'hfc78;
assign q[3695]= 16'h361;
assign q[3696]= 16'h9fe;
assign q[3697]= 16'h1029;
assign q[3698]= 16'h15bd;
assign q[3699]= 16'h1a98;
assign q[3700]= 16'h1e9d;
assign q[3701]= 16'h21b2;
assign q[3702]= 16'h23c2;
assign q[3703]= 16'h24bf;
assign q[3704]= 16'h24a4;
assign q[3705]= 16'h236f;
assign q[3706]= 16'h212a;
assign q[3707]= 16'h1de4;
assign q[3708]= 16'h19b6;
assign q[3709]= 16'h14bd;
assign q[3710]= 16'hf1f;
assign q[3711]= 16'h906;
assign q[3712]= 16'h29e;
assign q[3713]= 16'hfc1a;
assign q[3714]= 16'hf5aa;
assign q[3715]= 16'hef7f;
assign q[3716]= 16'he9c8;
assign q[3717]= 16'he4b0;
assign q[3718]= 16'he05d;
assign q[3719]= 16'hdcee;
assign q[3720]= 16'hda7a;
assign q[3721]= 16'hd912;
assign q[3722]= 16'hd8ba;
assign q[3723]= 16'hd96f;
assign q[3724]= 16'hdb25;
assign q[3725]= 16'hddc6;
assign q[3726]= 16'he137;
assign q[3727]= 16'he551;
assign q[3728]= 16'he9ee;
assign q[3729]= 16'heede;
assign q[3730]= 16'hf3f3;
assign q[3731]= 16'hf8fc;
assign q[3732]= 16'hfdcc;
assign q[3733]= 16'h236;
assign q[3734]= 16'h616;
assign q[3735]= 16'h94b;
assign q[3736]= 16'hbbb;
assign q[3737]= 16'hd58;
assign q[3738]= 16'he1a;
assign q[3739]= 16'he04;
assign q[3740]= 16'hd1f;
assign q[3741]= 16'hb81;
assign q[3742]= 16'h944;
assign q[3743]= 16'h68a;
assign q[3744]= 16'h37b;
assign q[3745]= 16'h41;
assign q[3746]= 16'hfd0a;
assign q[3747]= 16'hf9ff;
assign q[3748]= 16'hf74b;
assign q[3749]= 16'hf516;
assign q[3750]= 16'hf381;
assign q[3751]= 16'hf2a5;
assign q[3752]= 16'hf298;
assign q[3753]= 16'hf361;
assign q[3754]= 16'hf504;
assign q[3755]= 16'hf779;
assign q[3756]= 16'hfaaf;
assign q[3757]= 16'hfe8e;
assign q[3758]= 16'h2f5;
assign q[3759]= 16'h7c1;
assign q[3760]= 16'hcc6;
assign q[3761]= 16'h11d8;
assign q[3762]= 16'h16ca;
assign q[3763]= 16'h1b6d;
assign q[3764]= 16'h1f98;
assign q[3765]= 16'h2325;
assign q[3766]= 16'h25f1;
assign q[3767]= 16'h27e5;
assign q[3768]= 16'h28ed;
assign q[3769]= 16'h2902;
assign q[3770]= 16'h2821;
assign q[3771]= 16'h2655;
assign q[3772]= 16'h23af;
assign q[3773]= 16'h2047;
assign q[3774]= 16'h1c3e;
assign q[3775]= 16'h17b9;
assign q[3776]= 16'h12e3;
assign q[3777]= 16'hde9;
assign q[3778]= 16'h8f9;
assign q[3779]= 16'h440;
assign q[3780]= 16'hffea;
assign q[3781]= 16'hfc1c;
assign q[3782]= 16'hf8fa;
assign q[3783]= 16'hf69e;
assign q[3784]= 16'hf51f;
assign q[3785]= 16'hf487;
assign q[3786]= 16'hf4dc;
assign q[3787]= 16'hf61a;
assign q[3788]= 16'hf834;
assign q[3789]= 16'hfb18;
assign q[3790]= 16'hfeac;
assign q[3791]= 16'h2cf;
assign q[3792]= 16'h75f;
assign q[3793]= 16'hc36;
assign q[3794]= 16'h112b;
assign q[3795]= 16'h1617;
assign q[3796]= 16'h1ad2;
assign q[3797]= 16'h1f38;
assign q[3798]= 16'h232a;
assign q[3799]= 16'h268c;
assign q[3800]= 16'h2949;
assign q[3801]= 16'h2b51;
assign q[3802]= 16'h2c9d;
assign q[3803]= 16'h2d29;
assign q[3804]= 16'h2cfb;
assign q[3805]= 16'h2c1d;
assign q[3806]= 16'h2a9d;
assign q[3807]= 16'h2892;
assign q[3808]= 16'h2610;
assign q[3809]= 16'h2334;
assign q[3810]= 16'h2018;
assign q[3811]= 16'h1cd7;
assign q[3812]= 16'h198b;
assign q[3813]= 16'h164d;
assign q[3814]= 16'h1332;
assign q[3815]= 16'h104a;
assign q[3816]= 16'hda4;
assign q[3817]= 16'hb47;
assign q[3818]= 16'h937;
assign q[3819]= 16'h772;
assign q[3820]= 16'h5f3;
assign q[3821]= 16'h4af;
assign q[3822]= 16'h39a;
assign q[3823]= 16'h2a3;
assign q[3824]= 16'h1b8;
assign q[3825]= 16'hc7;
assign q[3826]= 16'hffbe;
assign q[3827]= 16'hfe8a;
assign q[3828]= 16'hfd1d;
assign q[3829]= 16'hfb6c;
assign q[3830]= 16'hf96d;
assign q[3831]= 16'hf71c;
assign q[3832]= 16'hf47b;
assign q[3833]= 16'hf18e;
assign q[3834]= 16'hee60;
assign q[3835]= 16'heaff;
assign q[3836]= 16'he77e;
assign q[3837]= 16'he3f4;
assign q[3838]= 16'he07a;
assign q[3839]= 16'hdd2a;
assign q[3840]= 16'hda22;
assign q[3841]= 16'hd77c;
assign q[3842]= 16'hd553;
assign q[3843]= 16'hd3bf;
assign q[3844]= 16'hd2d6;
assign q[3845]= 16'hd2a8;
assign q[3846]= 16'hd341;
assign q[3847]= 16'hd4a8;
assign q[3848]= 16'hd6de;
assign q[3849]= 16'hd9df;
assign q[3850]= 16'hdd9e;
assign q[3851]= 16'he20b;
assign q[3852]= 16'he711;
assign q[3853]= 16'hec95;
assign q[3854]= 16'hf27a;
assign q[3855]= 16'hf89e;
assign q[3856]= 16'hfedf;
assign q[3857]= 16'h518;
assign q[3858]= 16'hb29;
assign q[3859]= 16'h10f0;
assign q[3860]= 16'h164d;
assign q[3861]= 16'h1b26;
assign q[3862]= 16'h1f63;
assign q[3863]= 16'h22f3;
assign q[3864]= 16'h25c9;
assign q[3865]= 16'h27df;
assign q[3866]= 16'h2933;
assign q[3867]= 16'h29cb;
assign q[3868]= 16'h29b1;
assign q[3869]= 16'h28f4;
assign q[3870]= 16'h27a7;
assign q[3871]= 16'h25e3;
assign q[3872]= 16'h23c0;
assign q[3873]= 16'h215b;
assign q[3874]= 16'h1ed0;
assign q[3875]= 16'h1c3a;
assign q[3876]= 16'h19b7;
assign q[3877]= 16'h175e;
assign q[3878]= 16'h1546;
assign q[3879]= 16'h1383;
assign q[3880]= 16'h1225;
assign q[3881]= 16'h1137;
assign q[3882]= 16'h10bf;
assign q[3883]= 16'h10c1;
assign q[3884]= 16'h113b;
assign q[3885]= 16'h1227;
assign q[3886]= 16'h137c;
assign q[3887]= 16'h152d;
assign q[3888]= 16'h172b;
assign q[3889]= 16'h1963;
assign q[3890]= 16'h1bc3;
assign q[3891]= 16'h1e37;
assign q[3892]= 16'h20aa;
assign q[3893]= 16'h2309;
assign q[3894]= 16'h2541;
assign q[3895]= 16'h2741;
assign q[3896]= 16'h28f8;
assign q[3897]= 16'h2a59;
assign q[3898]= 16'h2b59;
assign q[3899]= 16'h2bf0;
assign q[3900]= 16'h2c16;
assign q[3901]= 16'h2bca;
assign q[3902]= 16'h2b09;
assign q[3903]= 16'h29d6;
assign q[3904]= 16'h2836;
assign q[3905]= 16'h262d;
assign q[3906]= 16'h23c5;
assign q[3907]= 16'h2106;
assign q[3908]= 16'h1dfd;
assign q[3909]= 16'h1ab6;
assign q[3910]= 16'h173e;
assign q[3911]= 16'h13a3;
assign q[3912]= 16'hff5;
assign q[3913]= 16'hc43;
assign q[3914]= 16'h89c;
assign q[3915]= 16'h50f;
assign q[3916]= 16'h1aa;
assign q[3917]= 16'hfe7f;
assign q[3918]= 16'hfb97;
assign q[3919]= 16'hf902;
assign q[3920]= 16'hf6ca;
assign q[3921]= 16'hf4fa;
assign q[3922]= 16'hf39b;
assign q[3923]= 16'hf2b4;
assign q[3924]= 16'hf24a;
assign q[3925]= 16'hf260;
assign q[3926]= 16'hf2f7;
assign q[3927]= 16'hf40e;
assign q[3928]= 16'hf59f;
assign q[3929]= 16'hf7a5;
assign q[3930]= 16'hfa17;
assign q[3931]= 16'hfce9;
assign q[3932]= 16'he;
assign q[3933]= 16'h377;
assign q[3934]= 16'h712;
assign q[3935]= 16'hacd;
assign q[3936]= 16'he93;
assign q[3937]= 16'h1252;
assign q[3938]= 16'h15f3;
assign q[3939]= 16'h1962;
assign q[3940]= 16'h1c8d;
assign q[3941]= 16'h1f5f;
assign q[3942]= 16'h21c9;
assign q[3943]= 16'h23ba;
assign q[3944]= 16'h2526;
assign q[3945]= 16'h2602;
assign q[3946]= 16'h2647;
assign q[3947]= 16'h25ef;
assign q[3948]= 16'h24fa;
assign q[3949]= 16'h2368;
assign q[3950]= 16'h213e;
assign q[3951]= 16'h1e83;
assign q[3952]= 16'h1b40;
assign q[3953]= 16'h1782;
assign q[3954]= 16'h1359;
assign q[3955]= 16'hed3;
assign q[3956]= 16'ha03;
assign q[3957]= 16'h4fc;
assign q[3958]= 16'hffd4;
assign q[3959]= 16'hfa9d;
assign q[3960]= 16'hf56c;
assign q[3961]= 16'hf056;
assign q[3962]= 16'heb6f;
assign q[3963]= 16'he6c9;
assign q[3964]= 16'he277;
assign q[3965]= 16'hde88;
assign q[3966]= 16'hdb0c;
assign q[3967]= 16'hd80f;
assign q[3968]= 16'hd59c;
assign q[3969]= 16'hd3bb;
assign q[3970]= 16'hd273;
assign q[3971]= 16'hd1c6;
assign q[3972]= 16'hd1b6;
assign q[3973]= 16'hd240;
assign q[3974]= 16'hd362;
assign q[3975]= 16'hd512;
assign q[3976]= 16'hd748;
assign q[3977]= 16'hd9f7;
assign q[3978]= 16'hdd11;
assign q[3979]= 16'he084;
assign q[3980]= 16'he43f;
assign q[3981]= 16'he82d;
assign q[3982]= 16'hec38;
assign q[3983]= 16'hf049;
assign q[3984]= 16'hf44a;
assign q[3985]= 16'hf825;
assign q[3986]= 16'hfbc2;
assign q[3987]= 16'hff0d;
assign q[3988]= 16'h1f0;
assign q[3989]= 16'h45d;
assign q[3990]= 16'h643;
assign q[3991]= 16'h797;
assign q[3992]= 16'h84e;
assign q[3993]= 16'h865;
assign q[3994]= 16'h7d8;
assign q[3995]= 16'h6ac;
assign q[3996]= 16'h4e5;
assign q[3997]= 16'h28d;
assign q[3998]= 16'hffb3;
assign q[3999]= 16'hfc64;
assign q[4000]= 16'hf8b4;
assign q[4001]= 16'hf4b9;
assign q[4002]= 16'hf088;
assign q[4003]= 16'hec39;
assign q[4004]= 16'he7e3;
assign q[4005]= 16'he39f;
assign q[4006]= 16'hdf81;
assign q[4007]= 16'hdb9f;
assign q[4008]= 16'hd80a;
assign q[4009]= 16'hd4d2;
assign q[4010]= 16'hd205;
assign q[4011]= 16'hcfab;
assign q[4012]= 16'hcdc9;
assign q[4013]= 16'hcc64;
assign q[4014]= 16'hcb78;
assign q[4015]= 16'hcb04;
assign q[4016]= 16'hcaff;
assign q[4017]= 16'hcb61;
assign q[4018]= 16'hcc1e;
assign q[4019]= 16'hcd29;
assign q[4020]= 16'hce75;
assign q[4021]= 16'hcff5;
assign q[4022]= 16'hd19a;
assign q[4023]= 16'hd358;
assign q[4024]= 16'hd523;
assign q[4025]= 16'hd6f1;
assign q[4026]= 16'hd8bb;
assign q[4027]= 16'hda79;
assign q[4028]= 16'hdc28;
assign q[4029]= 16'hddc6;
assign q[4030]= 16'hdf54;
assign q[4031]= 16'he0d3;
assign q[4032]= 16'he248;
assign q[4033]= 16'he3b7;
assign q[4034]= 16'he525;
assign q[4035]= 16'he69a;
assign q[4036]= 16'he81b;
assign q[4037]= 16'he9ad;
assign q[4038]= 16'heb56;
assign q[4039]= 16'hed1a;
assign q[4040]= 16'heef9;
assign q[4041]= 16'hf0f7;
assign q[4042]= 16'hf310;
assign q[4043]= 16'hf543;
assign q[4044]= 16'hf78a;
assign q[4045]= 16'hf9e0;
assign q[4046]= 16'hfc3d;
assign q[4047]= 16'hfe99;
assign q[4048]= 16'hea;
assign q[4049]= 16'h327;
assign q[4050]= 16'h548;
assign q[4051]= 16'h742;
assign q[4052]= 16'h90e;
assign q[4053]= 16'haa5;
assign q[4054]= 16'hc02;
assign q[4055]= 16'hd21;
assign q[4056]= 16'he01;
assign q[4057]= 16'hea3;
assign q[4058]= 16'hf08;
assign q[4059]= 16'hf37;
assign q[4060]= 16'hf36;
assign q[4061]= 16'hf0d;
assign q[4062]= 16'hec5;
assign q[4063]= 16'he6b;
assign q[4064]= 16'he09;
assign q[4065]= 16'hdab;
assign q[4066]= 16'hd5e;
assign q[4067]= 16'hd2b;
assign q[4068]= 16'hd1e;
assign q[4069]= 16'hd3f;
assign q[4070]= 16'hd96;
assign q[4071]= 16'he27;
assign q[4072]= 16'hef6;
assign q[4073]= 16'h1004;
assign q[4074]= 16'h114f;
assign q[4075]= 16'h12d5;
assign q[4076]= 16'h148f;
assign q[4077]= 16'h1676;
assign q[4078]= 16'h1881;
assign q[4079]= 16'h1aa6;
assign q[4080]= 16'h1cd8;
assign q[4081]= 16'h1f0e;
assign q[4082]= 16'h213a;
assign q[4083]= 16'h2350;
assign q[4084]= 16'h2547;
assign q[4085]= 16'h2714;
assign q[4086]= 16'h28ae;
assign q[4087]= 16'h2a10;
assign q[4088]= 16'h2b36;
assign q[4089]= 16'h2c1b;
assign q[4090]= 16'h2cc2;
assign q[4091]= 16'h2d2c;
assign q[4092]= 16'h2d5d;
assign q[4093]= 16'h2d5b;
assign q[4094]= 16'h2d30;
assign q[4095]= 16'h2ce5;
assign q[4096]= 16'h2c83;
assign q[4097]= 16'h2c17;
assign q[4098]= 16'h2bab;
assign q[4099]= 16'h2b4b;
assign q[4100]= 16'h2b01;
assign q[4101]= 16'h2ad4;
assign q[4102]= 16'h2acd;
assign q[4103]= 16'h2aef;
assign q[4104]= 16'h2b3d;
assign q[4105]= 16'h2bb6;
assign q[4106]= 16'h2c58;
assign q[4107]= 16'h2d1c;
assign q[4108]= 16'h2df9;
assign q[4109]= 16'h2ee4;
assign q[4110]= 16'h2fd0;
assign q[4111]= 16'h30ad;
assign q[4112]= 16'h316b;
assign q[4113]= 16'h31fa;
assign q[4114]= 16'h3248;
assign q[4115]= 16'h3245;
assign q[4116]= 16'h31e4;
assign q[4117]= 16'h3118;
assign q[4118]= 16'h2fd6;
assign q[4119]= 16'h2e1a;
assign q[4120]= 16'h2be1;
assign q[4121]= 16'h292b;
assign q[4122]= 16'h2601;
assign q[4123]= 16'h226b;
assign q[4124]= 16'h1e78;
assign q[4125]= 16'h1a3c;
assign q[4126]= 16'h15cb;
assign q[4127]= 16'h113f;
assign q[4128]= 16'hcb2;
assign q[4129]= 16'h840;
assign q[4130]= 16'h405;
assign q[4131]= 16'h1c;
assign q[4132]= 16'hfc9f;
assign q[4133]= 16'hf9a4;
assign q[4134]= 16'hf73d;
assign q[4135]= 16'hf57a;
assign q[4136]= 16'hf462;
assign q[4137]= 16'hf3f9;
assign q[4138]= 16'hf43d;
assign q[4139]= 16'hf523;
assign q[4140]= 16'hf69e;
assign q[4141]= 16'hf899;
assign q[4142]= 16'hfafa;
assign q[4143]= 16'hfda3;
assign q[4144]= 16'h72;
assign q[4145]= 16'h348;
assign q[4146]= 16'h5fe;
assign q[4147]= 16'h872;
assign q[4148]= 16'ha82;
assign q[4149]= 16'hc11;
assign q[4150]= 16'hd06;
assign q[4151]= 16'hd4c;
assign q[4152]= 16'hcd5;
assign q[4153]= 16'hb9c;
assign q[4154]= 16'h9a1;
assign q[4155]= 16'h6ec;
assign q[4156]= 16'h38e;
assign q[4157]= 16'hff9f;
assign q[4158]= 16'hfb3a;
assign q[4159]= 16'hf682;
assign q[4160]= 16'hf19e;
assign q[4161]= 16'hecb7;
assign q[4162]= 16'he7f7;
assign q[4163]= 16'he388;
assign q[4164]= 16'hdf92;
assign q[4165]= 16'hdc39;
assign q[4166]= 16'hd99c;
assign q[4167]= 16'hd7d3;
assign q[4168]= 16'hd6f1;
assign q[4169]= 16'hd6fe;
assign q[4170]= 16'hd7fc;
assign q[4171]= 16'hd9e2;
assign q[4172]= 16'hdca1;
assign q[4173]= 16'he020;
assign q[4174]= 16'he440;
assign q[4175]= 16'he8dc;
assign q[4176]= 16'hedcb;
assign q[4177]= 16'hf2e0;
assign q[4178]= 16'hf7ee;
assign q[4179]= 16'hfcc8;
assign q[4180]= 16'h142;
assign q[4181]= 16'h539;
assign q[4182]= 16'h889;
assign q[4183]= 16'hb19;
assign q[4184]= 16'hcd7;
assign q[4185]= 16'hdba;
assign q[4186]= 16'hdc1;
assign q[4187]= 16'hcf5;
assign q[4188]= 16'hb68;
assign q[4189]= 16'h933;
assign q[4190]= 16'h678;
assign q[4191]= 16'h35d;
assign q[4192]= 16'hd;
assign q[4193]= 16'hfcb5;
assign q[4194]= 16'hf983;
assign q[4195]= 16'hf6a4;
assign q[4196]= 16'hf440;
assign q[4197]= 16'hf27d;
assign q[4198]= 16'hf179;
assign q[4199]= 16'hf149;
assign q[4200]= 16'hf1fb;
assign q[4201]= 16'hf394;
assign q[4202]= 16'hf60c;
assign q[4203]= 16'hf956;
assign q[4204]= 16'hfd58;
assign q[4205]= 16'h1f1;
assign q[4206]= 16'h6f9;
assign q[4207]= 16'hc43;
assign q[4208]= 16'h119c;
assign q[4209]= 16'h16d2;
assign q[4210]= 16'h1bb0;
assign q[4211]= 16'h2004;
assign q[4212]= 16'h23a2;
assign q[4213]= 16'h2660;
assign q[4214]= 16'h281f;
assign q[4215]= 16'h28c5;
assign q[4216]= 16'h2846;
assign q[4217]= 16'h269e;
assign q[4218]= 16'h23d2;
assign q[4219]= 16'h1ff5;
assign q[4220]= 16'h1b22;
assign q[4221]= 16'h157d;
assign q[4222]= 16'hf32;
assign q[4223]= 16'h874;
assign q[4224]= 16'h17a;
assign q[4225]= 16'hfa7d;
assign q[4226]= 16'hf3b7;
assign q[4227]= 16'hed60;
assign q[4228]= 16'he7ad;
assign q[4229]= 16'he2cd;
assign q[4230]= 16'hdeea;
assign q[4231]= 16'hdc23;
assign q[4232]= 16'hda8e;
assign q[4233]= 16'hda39;
assign q[4234]= 16'hdb24;
assign q[4235]= 16'hdd48;
assign q[4236]= 16'he092;
assign q[4237]= 16'he4e7;
assign q[4238]= 16'hea22;
assign q[4239]= 16'hf018;
assign q[4240]= 16'hf69a;
assign q[4241]= 16'hfd75;
assign q[4242]= 16'h472;
assign q[4243]= 16'hb60;
assign q[4244]= 16'h120a;
assign q[4245]= 16'h1843;
assign q[4246]= 16'h1de1;
assign q[4247]= 16'h22c1;
assign q[4248]= 16'h26ca;
assign q[4249]= 16'h29e7;
assign q[4250]= 16'h2c10;
assign q[4251]= 16'h2d43;
assign q[4252]= 16'h2d87;
assign q[4253]= 16'h2cee;
assign q[4254]= 16'h2b8c;
assign q[4255]= 16'h2980;
assign q[4256]= 16'h26ea;
assign q[4257]= 16'h23ef;
assign q[4258]= 16'h20b6;
assign q[4259]= 16'h1d66;
assign q[4260]= 16'h1a26;
assign q[4261]= 16'h1718;
assign q[4262]= 16'h145d;
assign q[4263]= 16'h1211;
assign q[4264]= 16'h1048;
assign q[4265]= 16'hf12;
assign q[4266]= 16'he7a;
assign q[4267]= 16'he81;
assign q[4268]= 16'hf24;
assign q[4269]= 16'h105a;
assign q[4270]= 16'h1213;
assign q[4271]= 16'h143e;
assign q[4272]= 16'h16c3;
assign q[4273]= 16'h1989;
assign q[4274]= 16'h1c78;
assign q[4275]= 16'h1f73;
assign q[4276]= 16'h2263;
assign q[4277]= 16'h252f;
assign q[4278]= 16'h27c3;
assign q[4279]= 16'h2a0d;
assign q[4280]= 16'h2c00;
assign q[4281]= 16'h2d94;
assign q[4282]= 16'h2ec3;
assign q[4283]= 16'h2f8f;
assign q[4284]= 16'h2ffb;
assign q[4285]= 16'h3010;
assign q[4286]= 16'h2fda;
assign q[4287]= 16'h2f66;
assign q[4288]= 16'h2ec5;
assign q[4289]= 16'h2e09;
assign q[4290]= 16'h2d42;
assign q[4291]= 16'h2c82;
assign q[4292]= 16'h2bd8;
assign q[4293]= 16'h2b51;
assign q[4294]= 16'h2af8;
assign q[4295]= 16'h2ad4;
assign q[4296]= 16'h2aea;
assign q[4297]= 16'h2b39;
assign q[4298]= 16'h2bbe;
assign q[4299]= 16'h2c70;
assign q[4300]= 16'h2d47;
assign q[4301]= 16'h2e33;
assign q[4302]= 16'h2f25;
assign q[4303]= 16'h300a;
assign q[4304]= 16'h30d0;
assign q[4305]= 16'h3164;
assign q[4306]= 16'h31b1;
assign q[4307]= 16'h31a5;
assign q[4308]= 16'h3130;
assign q[4309]= 16'h3045;
assign q[4310]= 16'h2ed6;
assign q[4311]= 16'h2cde;
assign q[4312]= 16'h2a56;
assign q[4313]= 16'h2740;
assign q[4314]= 16'h239d;
assign q[4315]= 16'h1f75;
assign q[4316]= 16'h1ad3;
assign q[4317]= 16'h15c6;
assign q[4318]= 16'h105d;
assign q[4319]= 16'haac;
assign q[4320]= 16'h4c9;
assign q[4321]= 16'hfecc;
assign q[4322]= 16'hf8c8;
assign q[4323]= 16'hf2d6;
assign q[4324]= 16'hed0d;
assign q[4325]= 16'he782;
assign q[4326]= 16'he249;
assign q[4327]= 16'hdd72;
assign q[4328]= 16'hd90d;
assign q[4329]= 16'hd526;
assign q[4330]= 16'hd1c7;
assign q[4331]= 16'hcef4;
assign q[4332]= 16'hccb2;
assign q[4333]= 16'hcb01;
assign q[4334]= 16'hc9df;
assign q[4335]= 16'hc946;
assign q[4336]= 16'hc930;
assign q[4337]= 16'hc995;
assign q[4338]= 16'hca6a;
assign q[4339]= 16'hcba5;
assign q[4340]= 16'hcd3c;
assign q[4341]= 16'hcf22;
assign q[4342]= 16'hd14d;
assign q[4343]= 16'hd3b4;
assign q[4344]= 16'hd64c;
assign q[4345]= 16'hd90d;
assign q[4346]= 16'hdbf0;
assign q[4347]= 16'hdeef;
assign q[4348]= 16'he205;
assign q[4349]= 16'he52d;
assign q[4350]= 16'he864;
assign q[4351]= 16'heba8;
assign q[4352]= 16'heef7;
assign q[4353]= 16'hf24d;
assign q[4354]= 16'hf5a9;
assign q[4355]= 16'hf908;
assign q[4356]= 16'hfc65;
assign q[4357]= 16'hffbd;
assign q[4358]= 16'h309;
assign q[4359]= 16'h643;
assign q[4360]= 16'h963;
assign q[4361]= 16'hc60;
assign q[4362]= 16'hf2e;
assign q[4363]= 16'h11c4;
assign q[4364]= 16'h1416;
assign q[4365]= 16'h1616;
assign q[4366]= 16'h17bb;
assign q[4367]= 16'h18f7;
assign q[4368]= 16'h19c2;
assign q[4369]= 16'h1a11;
assign q[4370]= 16'h19df;
assign q[4371]= 16'h1926;
assign q[4372]= 16'h17e4;
assign q[4373]= 16'h161a;
assign q[4374]= 16'h13cb;
assign q[4375]= 16'h10ff;
assign q[4376]= 16'hdbf;
assign q[4377]= 16'ha19;
assign q[4378]= 16'h61c;
assign q[4379]= 16'h1dc;
assign q[4380]= 16'hfd6f;
assign q[4381]= 16'hf8e9;
assign q[4382]= 16'hf464;
assign q[4383]= 16'heff9;
assign q[4384]= 16'hebc1;
assign q[4385]= 16'he7d4;
assign q[4386]= 16'he449;
assign q[4387]= 16'he137;
assign q[4388]= 16'hdeb2;
assign q[4389]= 16'hdcc9;
assign q[4390]= 16'hdb8c;
assign q[4391]= 16'hdb03;
assign q[4392]= 16'hdb36;
assign q[4393]= 16'hdc28;
assign q[4394]= 16'hddd7;
assign q[4395]= 16'he040;
assign q[4396]= 16'he359;
assign q[4397]= 16'he716;
assign q[4398]= 16'heb6a;
assign q[4399]= 16'hf043;
assign q[4400]= 16'hf58c;
assign q[4401]= 16'hfb30;
assign q[4402]= 16'h118;
assign q[4403]= 16'h72c;
assign q[4404]= 16'hd55;
assign q[4405]= 16'h1378;
assign q[4406]= 16'h197f;
assign q[4407]= 16'h1f51;
assign q[4408]= 16'h24d9;
assign q[4409]= 16'h2a00;
assign q[4410]= 16'h2eb4;
assign q[4411]= 16'h32e3;
assign q[4412]= 16'h367d;
assign q[4413]= 16'h3974;
assign q[4414]= 16'h3bbe;
assign q[4415]= 16'h3d50;
assign q[4416]= 16'h3e25;
assign q[4417]= 16'h3e39;
assign q[4418]= 16'h3d8a;
assign q[4419]= 16'h3c19;
assign q[4420]= 16'h39eb;
assign q[4421]= 16'h3707;
assign q[4422]= 16'h3376;
assign q[4423]= 16'h2f45;
assign q[4424]= 16'h2a83;
assign q[4425]= 16'h2542;
assign q[4426]= 16'h1f96;
assign q[4427]= 16'h1995;
assign q[4428]= 16'h1358;
assign q[4429]= 16'hcf9;
assign q[4430]= 16'h693;
assign q[4431]= 16'h43;
assign q[4432]= 16'hfa24;
assign q[4433]= 16'hf451;
assign q[4434]= 16'heee6;
assign q[4435]= 16'he9fa;
assign q[4436]= 16'he5a6;
assign q[4437]= 16'he1fb;
assign q[4438]= 16'hdf0b;
assign q[4439]= 16'hdce2;
assign q[4440]= 16'hdb86;
assign q[4441]= 16'hdafb;
assign q[4442]= 16'hdb3f;
assign q[4443]= 16'hdc4a;
assign q[4444]= 16'hde12;
assign q[4445]= 16'he084;
assign q[4446]= 16'he38c;
assign q[4447]= 16'he712;
assign q[4448]= 16'heafa;
assign q[4449]= 16'hef27;
assign q[4450]= 16'hf378;
assign q[4451]= 16'hf7cf;
assign q[4452]= 16'hfc0c;
assign q[4453]= 16'h10;
assign q[4454]= 16'h3c2;
assign q[4455]= 16'h707;
assign q[4456]= 16'h9cb;
assign q[4457]= 16'hbfd;
assign q[4458]= 16'hd91;
assign q[4459]= 16'he81;
assign q[4460]= 16'heca;
assign q[4461]= 16'he6f;
assign q[4462]= 16'hd78;
assign q[4463]= 16'hbf2;
assign q[4464]= 16'h9eb;
assign q[4465]= 16'h776;
assign q[4466]= 16'h4a8;
assign q[4467]= 16'h197;
assign q[4468]= 16'hfe5b;
assign q[4469]= 16'hfb07;
assign q[4470]= 16'hf7b2;
assign q[4471]= 16'hf46e;
assign q[4472]= 16'hf14b;
assign q[4473]= 16'hee57;
assign q[4474]= 16'heb9c;
assign q[4475]= 16'he91f;
assign q[4476]= 16'he6e4;
assign q[4477]= 16'he4e9;
assign q[4478]= 16'he32c;
assign q[4479]= 16'he1a4;
assign q[4480]= 16'he04b;
assign q[4481]= 16'hdf14;
assign q[4482]= 16'hddf6;
assign q[4483]= 16'hdce6;
assign q[4484]= 16'hdbd9;
assign q[4485]= 16'hdac6;
assign q[4486]= 16'hd9a6;
assign q[4487]= 16'hd875;
assign q[4488]= 16'hd72f;
assign q[4489]= 16'hd5d8;
assign q[4490]= 16'hd471;
assign q[4491]= 16'hd303;
assign q[4492]= 16'hd198;
assign q[4493]= 16'hd03a;
assign q[4494]= 16'hcefa;
assign q[4495]= 16'hcde6;
assign q[4496]= 16'hcd0f;
assign q[4497]= 16'hcc84;
assign q[4498]= 16'hcc57;
assign q[4499]= 16'hcc95;
assign q[4500]= 16'hcd4b;
assign q[4501]= 16'hce84;
assign q[4502]= 16'hd045;
assign q[4503]= 16'hd295;
assign q[4504]= 16'hd572;
assign q[4505]= 16'hd8da;
assign q[4506]= 16'hdcc7;
assign q[4507]= 16'he12d;
assign q[4508]= 16'he601;
assign q[4509]= 16'heb32;
assign q[4510]= 16'hf0af;
assign q[4511]= 16'hf663;
assign q[4512]= 16'hfc3a;
assign q[4513]= 16'h21e;
assign q[4514]= 16'h7fc;
assign q[4515]= 16'hdbd;
assign q[4516]= 16'h134e;
assign q[4517]= 16'h189e;
assign q[4518]= 16'h1d9c;
assign q[4519]= 16'h223b;
assign q[4520]= 16'h266e;
assign q[4521]= 16'h2a2e;
assign q[4522]= 16'h2d72;
assign q[4523]= 16'h3037;
assign q[4524]= 16'h327b;
assign q[4525]= 16'h343e;
assign q[4526]= 16'h3581;
assign q[4527]= 16'h3647;
assign q[4528]= 16'h3695;
assign q[4529]= 16'h3671;
assign q[4530]= 16'h35df;
assign q[4531]= 16'h34e8;
assign q[4532]= 16'h3391;
assign q[4533]= 16'h31e1;
assign q[4534]= 16'h2fe1;
assign q[4535]= 16'h2d96;
assign q[4536]= 16'h2b08;
assign q[4537]= 16'h283d;
assign q[4538]= 16'h253c;
assign q[4539]= 16'h220d;
assign q[4540]= 16'h1eb5;
assign q[4541]= 16'h1b3c;
assign q[4542]= 16'h17a8;
assign q[4543]= 16'h1400;
assign q[4544]= 16'h104b;
assign q[4545]= 16'hc90;
assign q[4546]= 16'h8d5;
assign q[4547]= 16'h522;
assign q[4548]= 16'h17c;
assign q[4549]= 16'hfdeb;
assign q[4550]= 16'hfa71;
assign q[4551]= 16'hf716;
assign q[4552]= 16'hf3de;
assign q[4553]= 16'hf0cc;
assign q[4554]= 16'hede2;
assign q[4555]= 16'heb24;
assign q[4556]= 16'he891;
assign q[4557]= 16'he62c;
assign q[4558]= 16'he3f4;
assign q[4559]= 16'he1e8;
assign q[4560]= 16'he008;
assign q[4561]= 16'hde53;
assign q[4562]= 16'hdcc8;
assign q[4563]= 16'hdb65;
assign q[4564]= 16'hda2c;
assign q[4565]= 16'hd91b;
assign q[4566]= 16'hd834;
assign q[4567]= 16'hd778;
assign q[4568]= 16'hd6e9;
assign q[4569]= 16'hd68b;
assign q[4570]= 16'hd661;
assign q[4571]= 16'hd66f;
assign q[4572]= 16'hd6b9;
assign q[4573]= 16'hd745;
assign q[4574]= 16'hd817;
assign q[4575]= 16'hd934;
assign q[4576]= 16'hda9e;
assign q[4577]= 16'hdc59;
assign q[4578]= 16'hde66;
assign q[4579]= 16'he0c6;
assign q[4580]= 16'he377;
assign q[4581]= 16'he677;
assign q[4582]= 16'he9c1;
assign q[4583]= 16'hed4e;
assign q[4584]= 16'hf117;
assign q[4585]= 16'hf511;
assign q[4586]= 16'hf931;
assign q[4587]= 16'hfd6b;
assign q[4588]= 16'h1b1;
assign q[4589]= 16'h5f5;
assign q[4590]= 16'ha2a;
assign q[4591]= 16'he3f;
assign q[4592]= 16'h1226;
assign q[4593]= 16'h15d2;
assign q[4594]= 16'h1935;
assign q[4595]= 16'h1c44;
assign q[4596]= 16'h1ef3;
assign q[4597]= 16'h2139;
assign q[4598]= 16'h230d;
assign q[4599]= 16'h246a;
assign q[4600]= 16'h2549;
assign q[4601]= 16'h25a9;
assign q[4602]= 16'h2586;
assign q[4603]= 16'h24e0;
assign q[4604]= 16'h23b9;
assign q[4605]= 16'h2212;
assign q[4606]= 16'h1fee;
assign q[4607]= 16'h1d53;
assign q[4608]= 16'h1a47;
assign q[4609]= 16'h16d0;
assign q[4610]= 16'h12f8;
assign q[4611]= 16'hec7;
assign q[4612]= 16'ha49;
assign q[4613]= 16'h58a;
assign q[4614]= 16'h98;
assign q[4615]= 16'hfb84;
assign q[4616]= 16'hf65c;
assign q[4617]= 16'hf133;
assign q[4618]= 16'hec1d;
assign q[4619]= 16'he72d;
assign q[4620]= 16'he27a;
assign q[4621]= 16'hde17;
assign q[4622]= 16'hda1c;
assign q[4623]= 16'hd69d;
assign q[4624]= 16'hd3ad;
assign q[4625]= 16'hd161;
assign q[4626]= 16'hcfc8;
assign q[4627]= 16'hcef0;
assign q[4628]= 16'hcee4;
assign q[4629]= 16'hcfaa;
assign q[4630]= 16'hd144;
assign q[4631]= 16'hd3b1;
assign q[4632]= 16'hd6e8;
assign q[4633]= 16'hdade;
assign q[4634]= 16'hdf81;
assign q[4635]= 16'he4bc;
assign q[4636]= 16'hea73;
assign q[4637]= 16'hf088;
assign q[4638]= 16'hf6db;
assign q[4639]= 16'hfd46;
assign q[4640]= 16'h3a4;
assign q[4641]= 16'h9d2;
assign q[4642]= 16'hfa9;
assign q[4643]= 16'h1507;
assign q[4644]= 16'h19cc;
assign q[4645]= 16'h1ddb;
assign q[4646]= 16'h211d;
assign q[4647]= 16'h2382;
assign q[4648]= 16'h24fe;
assign q[4649]= 16'h258c;
assign q[4650]= 16'h252f;
assign q[4651]= 16'h23f2;
assign q[4652]= 16'h21e3;
assign q[4653]= 16'h1f19;
assign q[4654]= 16'h1bb1;
assign q[4655]= 16'h17cb;
assign q[4656]= 16'h138c;
assign q[4657]= 16'hf19;
assign q[4658]= 16'ha9c;
assign q[4659]= 16'h63c;
assign q[4660]= 16'h21f;
assign q[4661]= 16'hfe6b;
assign q[4662]= 16'hfb3e;
assign q[4663]= 16'hf8b5;
assign q[4664]= 16'hf6e5;
assign q[4665]= 16'hf5de;
assign q[4666]= 16'hf5a9;
assign q[4667]= 16'hf64a;
assign q[4668]= 16'hf7bb;
assign q[4669]= 16'hf9f2;
assign q[4670]= 16'hfcdd;
assign q[4671]= 16'h68;
assign q[4672]= 16'h478;
assign q[4673]= 16'h8ef;
assign q[4674]= 16'hdaf;
assign q[4675]= 16'h1295;
assign q[4676]= 16'h1782;
assign q[4677]= 16'h1c55;
assign q[4678]= 16'h20f1;
assign q[4679]= 16'h253c;
assign q[4680]= 16'h291f;
assign q[4681]= 16'h2c88;
assign q[4682]= 16'h2f6a;
assign q[4683]= 16'h31bd;
assign q[4684]= 16'h337d;
assign q[4685]= 16'h34ab;
assign q[4686]= 16'h354f;
assign q[4687]= 16'h3572;
assign q[4688]= 16'h3520;
assign q[4689]= 16'h346b;
assign q[4690]= 16'h3362;
assign q[4691]= 16'h3218;
assign q[4692]= 16'h309f;
assign q[4693]= 16'h2f08;
assign q[4694]= 16'h2d63;
assign q[4695]= 16'h2bbd;
assign q[4696]= 16'h2a21;
assign q[4697]= 16'h2897;
assign q[4698]= 16'h2723;
assign q[4699]= 16'h25c7;
assign q[4700]= 16'h2481;
assign q[4701]= 16'h234d;
assign q[4702]= 16'h2223;
assign q[4703]= 16'h20fa;
assign q[4704]= 16'h1fc9;
assign q[4705]= 16'h1e84;
assign q[4706]= 16'h1d1f;
assign q[4707]= 16'h1b8f;
assign q[4708]= 16'h19cb;
assign q[4709]= 16'h17ca;
assign q[4710]= 16'h1586;
assign q[4711]= 16'h12fa;
assign q[4712]= 16'h1025;
assign q[4713]= 16'hd09;
assign q[4714]= 16'h9a9;
assign q[4715]= 16'h60c;
assign q[4716]= 16'h23b;
assign q[4717]= 16'hfe42;
assign q[4718]= 16'hfa2b;
assign q[4719]= 16'hf606;
assign q[4720]= 16'hf1e1;
assign q[4721]= 16'hedcb;
assign q[4722]= 16'he9d2;
assign q[4723]= 16'he604;
assign q[4724]= 16'he26e;
assign q[4725]= 16'hdf19;
assign q[4726]= 16'hdc10;
assign q[4727]= 16'hd959;
assign q[4728]= 16'hd6f8;
assign q[4729]= 16'hd4f0;
assign q[4730]= 16'hd342;
assign q[4731]= 16'hd1ea;
assign q[4732]= 16'hd0e6;
assign q[4733]= 16'hd030;
assign q[4734]= 16'hcfc1;
assign q[4735]= 16'hcf91;
assign q[4736]= 16'hcf97;
assign q[4737]= 16'hcfcb;
assign q[4738]= 16'hd023;
assign q[4739]= 16'hd098;
assign q[4740]= 16'hd120;
assign q[4741]= 16'hd1b4;
assign q[4742]= 16'hd24d;
assign q[4743]= 16'hd2e5;
assign q[4744]= 16'hd377;
assign q[4745]= 16'hd3ff;
assign q[4746]= 16'hd47a;
assign q[4747]= 16'hd4e6;
assign q[4748]= 16'hd540;
assign q[4749]= 16'hd587;
assign q[4750]= 16'hd5bc;
assign q[4751]= 16'hd5dd;
assign q[4752]= 16'hd5ec;
assign q[4753]= 16'hd5e7;
assign q[4754]= 16'hd5d1;
assign q[4755]= 16'hd5a9;
assign q[4756]= 16'hd570;
assign q[4757]= 16'hd528;
assign q[4758]= 16'hd4d1;
assign q[4759]= 16'hd46e;
assign q[4760]= 16'hd3ff;
assign q[4761]= 16'hd388;
assign q[4762]= 16'hd30c;
assign q[4763]= 16'hd28e;
assign q[4764]= 16'hd212;
assign q[4765]= 16'hd19d;
assign q[4766]= 16'hd133;
assign q[4767]= 16'hd0db;
assign q[4768]= 16'hd099;
assign q[4769]= 16'hd075;
assign q[4770]= 16'hd074;
assign q[4771]= 16'hd09b;
assign q[4772]= 16'hd0ef;
assign q[4773]= 16'hd174;
assign q[4774]= 16'hd22e;
assign q[4775]= 16'hd31f;
assign q[4776]= 16'hd446;
assign q[4777]= 16'hd5a3;
assign q[4778]= 16'hd732;
assign q[4779]= 16'hd8ef;
assign q[4780]= 16'hdad4;
assign q[4781]= 16'hdcd9;
assign q[4782]= 16'hdef4;
assign q[4783]= 16'he119;
assign q[4784]= 16'he33f;
assign q[4785]= 16'he558;
assign q[4786]= 16'he758;
assign q[4787]= 16'he931;
assign q[4788]= 16'heada;
assign q[4789]= 16'hec45;
assign q[4790]= 16'hed6a;
assign q[4791]= 16'hee40;
assign q[4792]= 16'heec1;
assign q[4793]= 16'heee9;
assign q[4794]= 16'heeb7;
assign q[4795]= 16'hee2a;
assign q[4796]= 16'hed46;
assign q[4797]= 16'hec10;
assign q[4798]= 16'hea8f;
assign q[4799]= 16'he8cc;
assign q[4800]= 16'he6d3;
assign q[4801]= 16'he4ae;
assign q[4802]= 16'he26b;
assign q[4803]= 16'he016;
assign q[4804]= 16'hddbe;
assign q[4805]= 16'hdb6e;
assign q[4806]= 16'hd933;
assign q[4807]= 16'hd717;
assign q[4808]= 16'hd525;
assign q[4809]= 16'hd366;
assign q[4810]= 16'hd1de;
assign q[4811]= 16'hd095;
assign q[4812]= 16'hcf8d;
assign q[4813]= 16'hcec9;
assign q[4814]= 16'hce48;
assign q[4815]= 16'hce0b;
assign q[4816]= 16'hce10;
assign q[4817]= 16'hce54;
assign q[4818]= 16'hced6;
assign q[4819]= 16'hcf93;
assign q[4820]= 16'hd087;
assign q[4821]= 16'hd1b1;
assign q[4822]= 16'hd30f;
assign q[4823]= 16'hd49f;
assign q[4824]= 16'hd660;
assign q[4825]= 16'hd852;
assign q[4826]= 16'hda76;
assign q[4827]= 16'hdccb;
assign q[4828]= 16'hdf53;
assign q[4829]= 16'he20f;
assign q[4830]= 16'he4fe;
assign q[4831]= 16'he821;
assign q[4832]= 16'heb77;
assign q[4833]= 16'heefe;
assign q[4834]= 16'hf2b4;
assign q[4835]= 16'hf694;
assign q[4836]= 16'hfa97;
assign q[4837]= 16'hfeb8;
assign q[4838]= 16'h2ec;
assign q[4839]= 16'h72a;
assign q[4840]= 16'hb67;
assign q[4841]= 16'hf95;
assign q[4842]= 16'h13a8;
assign q[4843]= 16'h1791;
assign q[4844]= 16'h1b43;
assign q[4845]= 16'h1eae;
assign q[4846]= 16'h21c6;
assign q[4847]= 16'h247d;
assign q[4848]= 16'h26c9;
assign q[4849]= 16'h289f;
assign q[4850]= 16'h29f6;
assign q[4851]= 16'h2ac7;
assign q[4852]= 16'h2b0e;
assign q[4853]= 16'h2ac8;
assign q[4854]= 16'h29f4;
assign q[4855]= 16'h2893;
assign q[4856]= 16'h26a8;
assign q[4857]= 16'h2438;
assign q[4858]= 16'h2149;
assign q[4859]= 16'h1de3;
assign q[4860]= 16'h1a10;
assign q[4861]= 16'h15d9;
assign q[4862]= 16'h1149;
assign q[4863]= 16'hc6d;
assign q[4864]= 16'h750;
assign q[4865]= 16'h200;
assign q[4866]= 16'hfc8c;
assign q[4867]= 16'hf6ff;
assign q[4868]= 16'hf168;
assign q[4869]= 16'hebd7;
assign q[4870]= 16'he65b;
assign q[4871]= 16'he104;
assign q[4872]= 16'hdbe1;
assign q[4873]= 16'hd704;
assign q[4874]= 16'hd27c;
assign q[4875]= 16'hce5c;
assign q[4876]= 16'hcab2;
assign q[4877]= 16'hc791;
assign q[4878]= 16'hc507;
assign q[4879]= 16'hc323;
assign q[4880]= 16'hc1f2;
assign q[4881]= 16'hc180;
assign q[4882]= 16'hc1d4;
assign q[4883]= 16'hc2f5;
assign q[4884]= 16'hc4e5;
assign q[4885]= 16'hc7a3;
assign q[4886]= 16'hcb2a;
assign q[4887]= 16'hcf70;
assign q[4888]= 16'hd466;
assign q[4889]= 16'hd9fa;
assign q[4890]= 16'he014;
assign q[4891]= 16'he69b;
assign q[4892]= 16'hed6d;
assign q[4893]= 16'hf46b;
assign q[4894]= 16'hfb6f;
assign q[4895]= 16'h252;
assign q[4896]= 16'h8ef;
assign q[4897]= 16'hf20;
assign q[4898]= 16'h14c1;
assign q[4899]= 16'h19ae;
assign q[4900]= 16'h1dca;
assign q[4901]= 16'h20fb;
assign q[4902]= 16'h232d;
assign q[4903]= 16'h2452;
assign q[4904]= 16'h2464;
assign q[4905]= 16'h2361;
assign q[4906]= 16'h2153;
assign q[4907]= 16'h1e49;
assign q[4908]= 16'h1a58;
assign q[4909]= 16'h159d;
assign q[4910]= 16'h103b;
assign q[4911]= 16'ha59;
assign q[4912]= 16'h422;
assign q[4913]= 16'hfdc4;
assign q[4914]= 16'hf76c;
assign q[4915]= 16'hf149;
assign q[4916]= 16'heb87;
assign q[4917]= 16'he64e;
assign q[4918]= 16'he1c4;
assign q[4919]= 16'hde06;
assign q[4920]= 16'hdb2e;
assign q[4921]= 16'hd94c;
assign q[4922]= 16'hd86a;
assign q[4923]= 16'hd889;
assign q[4924]= 16'hd9a3;
assign q[4925]= 16'hdba8;
assign q[4926]= 16'hde85;
assign q[4927]= 16'he21d;
assign q[4928]= 16'he650;
assign q[4929]= 16'heafa;
assign q[4930]= 16'heff3;
assign q[4931]= 16'hf515;
assign q[4932]= 16'hfa36;
assign q[4933]= 16'hff31;
assign q[4934]= 16'h3e2;
assign q[4935]= 16'h82c;
assign q[4936]= 16'hbf5;
assign q[4937]= 16'hf29;
assign q[4938]= 16'h11bb;
assign q[4939]= 16'h13a6;
assign q[4940]= 16'h14eb;
assign q[4941]= 16'h1592;
assign q[4942]= 16'h15a9;
assign q[4943]= 16'h1543;
assign q[4944]= 16'h1479;
assign q[4945]= 16'h1366;
assign q[4946]= 16'h1227;
assign q[4947]= 16'h10dc;
assign q[4948]= 16'hfa3;
assign q[4949]= 16'he97;
assign q[4950]= 16'hdd2;
assign q[4951]= 16'hd69;
assign q[4952]= 16'hd6d;
assign q[4953]= 16'hde7;
assign q[4954]= 16'hede;
assign q[4955]= 16'h104f;
assign q[4956]= 16'h1232;
assign q[4957]= 16'h147b;
assign q[4958]= 16'h1716;
assign q[4959]= 16'h19ec;
assign q[4960]= 16'h1ce4;
assign q[4961]= 16'h1fe0;
assign q[4962]= 16'h22c3;
assign q[4963]= 16'h2571;
assign q[4964]= 16'h27cd;
assign q[4965]= 16'h29bf;
assign q[4966]= 16'h2b32;
assign q[4967]= 16'h2c18;
assign q[4968]= 16'h2c65;
assign q[4969]= 16'h2c16;
assign q[4970]= 16'h2b2d;
assign q[4971]= 16'h29b4;
assign q[4972]= 16'h27b8;
assign q[4973]= 16'h2550;
assign q[4974]= 16'h2293;
assign q[4975]= 16'h1f9f;
assign q[4976]= 16'h1c94;
assign q[4977]= 16'h1991;
assign q[4978]= 16'h16b9;
assign q[4979]= 16'h142a;
assign q[4980]= 16'h1201;
assign q[4981]= 16'h1057;
assign q[4982]= 16'hf3e;
assign q[4983]= 16'hec4;
assign q[4984]= 16'hef0;
assign q[4985]= 16'hfc2;
assign q[4986]= 16'h1131;
assign q[4987]= 16'h1330;
assign q[4988]= 16'h15aa;
assign q[4989]= 16'h1882;
assign q[4990]= 16'h1b9b;
assign q[4991]= 16'h1ed0;
assign q[4992]= 16'h21fb;
assign q[4993]= 16'h24f5;
assign q[4994]= 16'h2798;
assign q[4995]= 16'h29c0;
assign q[4996]= 16'h2b4c;
assign q[4997]= 16'h2c1f;
assign q[4998]= 16'h2c24;
assign q[4999]= 16'h2b4b;
assign q[5000]= 16'h298b;
assign q[5001]= 16'h26e5;
assign q[5002]= 16'h2361;
assign q[5003]= 16'h1f0d;
assign q[5004]= 16'h1a02;
assign q[5005]= 16'h145b;
assign q[5006]= 16'he3c;
assign q[5007]= 16'h7cd;
assign q[5008]= 16'h137;
assign q[5009]= 16'hfaa7;
assign q[5010]= 16'hf447;
assign q[5011]= 16'hee42;
assign q[5012]= 16'he8c1;
assign q[5013]= 16'he3e6;
assign q[5014]= 16'hdfcf;
assign q[5015]= 16'hdc94;
assign q[5016]= 16'hda48;
assign q[5017]= 16'hd8f2;
assign q[5018]= 16'hd895;
assign q[5019]= 16'hd92c;
assign q[5020]= 16'hdaab;
assign q[5021]= 16'hdcfe;
assign q[5022]= 16'he00e;
assign q[5023]= 16'he3bd;
assign q[5024]= 16'he7eb;
assign q[5025]= 16'hec76;
assign q[5026]= 16'hf139;
assign q[5027]= 16'hf611;
assign q[5028]= 16'hfadd;
assign q[5029]= 16'hff7c;
assign q[5030]= 16'h3d2;
assign q[5031]= 16'h7ca;
assign q[5032]= 16'hb4f;
assign q[5033]= 16'he54;
assign q[5034]= 16'h10d0;
assign q[5035]= 16'h12c1;
assign q[5036]= 16'h1429;
assign q[5037]= 16'h150f;
assign q[5038]= 16'h157d;
assign q[5039]= 16'h1582;
assign q[5040]= 16'h152f;
assign q[5041]= 16'h1495;
assign q[5042]= 16'h13c8;
assign q[5043]= 16'h12db;
assign q[5044]= 16'h11e1;
assign q[5045]= 16'h10e9;
assign q[5046]= 16'h1002;
assign q[5047]= 16'hf38;
assign q[5048]= 16'he94;
assign q[5049]= 16'he1b;
assign q[5050]= 16'hdcf;
assign q[5051]= 16'hdaf;
assign q[5052]= 16'hdb9;
assign q[5053]= 16'hde5;
assign q[5054]= 16'he2a;
assign q[5055]= 16'he7e;
assign q[5056]= 16'hed6;
assign q[5057]= 16'hf25;
assign q[5058]= 16'hf5e;
assign q[5059]= 16'hf76;
assign q[5060]= 16'hf60;
assign q[5061]= 16'hf12;
assign q[5062]= 16'he83;
assign q[5063]= 16'hdac;
assign q[5064]= 16'hc87;
assign q[5065]= 16'hb10;
assign q[5066]= 16'h946;
assign q[5067]= 16'h728;
assign q[5068]= 16'h4b9;
assign q[5069]= 16'h1fb;
assign q[5070]= 16'hfef6;
assign q[5071]= 16'hfbae;
assign q[5072]= 16'hf82a;
assign q[5073]= 16'hf475;
assign q[5074]= 16'hf098;
assign q[5075]= 16'hec9d;
assign q[5076]= 16'he88f;
assign q[5077]= 16'he47c;
assign q[5078]= 16'he06f;
assign q[5079]= 16'hdc75;
assign q[5080]= 16'hd89c;
assign q[5081]= 16'hd4f2;
assign q[5082]= 16'hd186;
assign q[5083]= 16'hce66;
assign q[5084]= 16'hcba0;
assign q[5085]= 16'hc943;
assign q[5086]= 16'hc75c;
assign q[5087]= 16'hc5f9;
assign q[5088]= 16'hc525;
assign q[5089]= 16'hc4eb;
assign q[5090]= 16'hc554;
assign q[5091]= 16'hc666;
assign q[5092]= 16'hc825;
assign q[5093]= 16'hca91;
assign q[5094]= 16'hcda8;
assign q[5095]= 16'hd164;
assign q[5096]= 16'hd5bc;
assign q[5097]= 16'hdaa0;
assign q[5098]= 16'he001;
assign q[5099]= 16'he5ca;
assign q[5100]= 16'hebe2;
assign q[5101]= 16'hf22f;
assign q[5102]= 16'hf893;
assign q[5103]= 16'hfeef;
assign q[5104]= 16'h523;
assign q[5105]= 16'hb0f;
assign q[5106]= 16'h1093;
assign q[5107]= 16'h1592;
assign q[5108]= 16'h19ee;
assign q[5109]= 16'h1d8f;
assign q[5110]= 16'h205f;
assign q[5111]= 16'h224f;
assign q[5112]= 16'h2351;
assign q[5113]= 16'h235f;
assign q[5114]= 16'h2279;
assign q[5115]= 16'h20a2;
assign q[5116]= 16'h1de5;
assign q[5117]= 16'h1a51;
assign q[5118]= 16'h15fa;
assign q[5119]= 16'h10f9;
assign q[5120]= 16'hb69;
assign q[5121]= 16'h56a;
assign q[5122]= 16'hff1e;
assign q[5123]= 16'hf8a4;
assign q[5124]= 16'hf21f;
assign q[5125]= 16'hebb2;
assign q[5126]= 16'he57b;
assign q[5127]= 16'hdf98;
assign q[5128]= 16'hda24;
assign q[5129]= 16'hd536;
assign q[5130]= 16'hd0e0;
assign q[5131]= 16'hcd30;
assign q[5132]= 16'hca32;
assign q[5133]= 16'hc7e9;
assign q[5134]= 16'hc658;
assign q[5135]= 16'hc57c;
assign q[5136]= 16'hc54d;
assign q[5137]= 16'hc5c3;
assign q[5138]= 16'hc6d0;
assign q[5139]= 16'hc865;
assign q[5140]= 16'hca74;
assign q[5141]= 16'hcceb;
assign q[5142]= 16'hcfb8;
assign q[5143]= 16'hd2cb;
assign q[5144]= 16'hd613;
assign q[5145]= 16'hd982;
assign q[5146]= 16'hdd09;
assign q[5147]= 16'he09e;
assign q[5148]= 16'he434;
assign q[5149]= 16'he7c5;
assign q[5150]= 16'heb4a;
assign q[5151]= 16'heebe;
assign q[5152]= 16'hf21c;
assign q[5153]= 16'hf563;
assign q[5154]= 16'hf892;
assign q[5155]= 16'hfba6;
assign q[5156]= 16'hfe9f;
assign q[5157]= 16'h17c;
assign q[5158]= 16'h43c;
assign q[5159]= 16'h6dd;
assign q[5160]= 16'h95c;
assign q[5161]= 16'hbb5;
assign q[5162]= 16'hde5;
assign q[5163]= 16'hfe5;
assign q[5164]= 16'h11b1;
assign q[5165]= 16'h1340;
assign q[5166]= 16'h148c;
assign q[5167]= 16'h158e;
assign q[5168]= 16'h163f;
assign q[5169]= 16'h1699;
assign q[5170]= 16'h1694;
assign q[5171]= 16'h162e;
assign q[5172]= 16'h1563;
assign q[5173]= 16'h1430;
assign q[5174]= 16'h1297;
assign q[5175]= 16'h1099;
assign q[5176]= 16'he3a;
assign q[5177]= 16'hb81;
assign q[5178]= 16'h874;
assign q[5179]= 16'h51f;
assign q[5180]= 16'h18c;
assign q[5181]= 16'hfdca;
assign q[5182]= 16'hf9e3;
assign q[5183]= 16'hf5e7;
assign q[5184]= 16'hf1e5;
assign q[5185]= 16'hedeb;
assign q[5186]= 16'hea08;
assign q[5187]= 16'he649;
assign q[5188]= 16'he2bb;
assign q[5189]= 16'hdf67;
assign q[5190]= 16'hdc57;
assign q[5191]= 16'hd993;
assign q[5192]= 16'hd720;
assign q[5193]= 16'hd501;
assign q[5194]= 16'hd338;
assign q[5195]= 16'hd1c5;
assign q[5196]= 16'hd0a6;
assign q[5197]= 16'hcfd6;
assign q[5198]= 16'hcf51;
assign q[5199]= 16'hcf12;
assign q[5200]= 16'hcf11;
assign q[5201]= 16'hcf48;
assign q[5202]= 16'hcfb0;
assign q[5203]= 16'hd041;
assign q[5204]= 16'hd0f6;
assign q[5205]= 16'hd1c9;
assign q[5206]= 16'hd2b4;
assign q[5207]= 16'hd3b4;
assign q[5208]= 16'hd4c6;
assign q[5209]= 16'hd5e9;
assign q[5210]= 16'hd71a;
assign q[5211]= 16'hd85b;
assign q[5212]= 16'hd9ab;
assign q[5213]= 16'hdb0d;
assign q[5214]= 16'hdc82;
assign q[5215]= 16'hde0d;
assign q[5216]= 16'hdfae;
assign q[5217]= 16'he167;
assign q[5218]= 16'he33a;
assign q[5219]= 16'he527;
assign q[5220]= 16'he72e;
assign q[5221]= 16'he94e;
assign q[5222]= 16'heb83;
assign q[5223]= 16'hedcd;
assign q[5224]= 16'hf025;
assign q[5225]= 16'hf288;
assign q[5226]= 16'hf4f0;
assign q[5227]= 16'hf757;
assign q[5228]= 16'hf9b6;
assign q[5229]= 16'hfc06;
assign q[5230]= 16'hfe41;
assign q[5231]= 16'h5f;
assign q[5232]= 16'h25c;
assign q[5233]= 16'h430;
assign q[5234]= 16'h5d8;
assign q[5235]= 16'h74e;
assign q[5236]= 16'h88f;
assign q[5237]= 16'h998;
assign q[5238]= 16'ha67;
assign q[5239]= 16'hafa;
assign q[5240]= 16'hb51;
assign q[5241]= 16'hb6c;
assign q[5242]= 16'hb4a;
assign q[5243]= 16'haee;
assign q[5244]= 16'ha57;
assign q[5245]= 16'h987;
assign q[5246]= 16'h87f;
assign q[5247]= 16'h741;
assign q[5248]= 16'h5cd;
assign q[5249]= 16'h425;
assign q[5250]= 16'h24b;
assign q[5251]= 16'h41;
assign q[5252]= 16'hfe0a;
assign q[5253]= 16'hfba7;
assign q[5254]= 16'hf91d;
assign q[5255]= 16'hf670;
assign q[5256]= 16'hf3a6;
assign q[5257]= 16'hf0c4;
assign q[5258]= 16'hedd4;
assign q[5259]= 16'headd;
assign q[5260]= 16'he7e8;
assign q[5261]= 16'he502;
assign q[5262]= 16'he234;
assign q[5263]= 16'hdf8c;
assign q[5264]= 16'hdd15;
assign q[5265]= 16'hdadb;
assign q[5266]= 16'hd8ea;
assign q[5267]= 16'hd74c;
assign q[5268]= 16'hd60a;
assign q[5269]= 16'hd52b;
assign q[5270]= 16'hd4b5;
assign q[5271]= 16'hd4aa;
assign q[5272]= 16'hd50b;
assign q[5273]= 16'hd5d3;
assign q[5274]= 16'hd6fe;
assign q[5275]= 16'hd882;
assign q[5276]= 16'hda54;
assign q[5277]= 16'hdc65;
assign q[5278]= 16'hdea6;
assign q[5279]= 16'he106;
assign q[5280]= 16'he371;
assign q[5281]= 16'he5d4;
assign q[5282]= 16'he81f;
assign q[5283]= 16'hea3e;
assign q[5284]= 16'hec24;
assign q[5285]= 16'hedc2;
assign q[5286]= 16'hef0f;
assign q[5287]= 16'hf005;
assign q[5288]= 16'hf0a1;
assign q[5289]= 16'hf0e4;
assign q[5290]= 16'hf0d5;
assign q[5291]= 16'hf07b;
assign q[5292]= 16'hefe6;
assign q[5293]= 16'hef24;
assign q[5294]= 16'hee4a;
assign q[5295]= 16'hed6d;
assign q[5296]= 16'heca2;
assign q[5297]= 16'hec00;
assign q[5298]= 16'heb9d;
assign q[5299]= 16'heb8e;
assign q[5300]= 16'hebe3;
assign q[5301]= 16'hecac;
assign q[5302]= 16'hedf4;
assign q[5303]= 16'hefc0;
assign q[5304]= 16'hf212;
assign q[5305]= 16'hf4e7;
assign q[5306]= 16'hf835;
assign q[5307]= 16'hfbee;
assign q[5308]= 16'h0;
assign q[5309]= 16'h455;
assign q[5310]= 16'h8d4;
assign q[5311]= 16'hd60;
assign q[5312]= 16'h11dc;
assign q[5313]= 16'h162a;
assign q[5314]= 16'h1a2c;
assign q[5315]= 16'h1dc5;
assign q[5316]= 16'h20de;
assign q[5317]= 16'h235f;
assign q[5318]= 16'h2538;
assign q[5319]= 16'h265a;
assign q[5320]= 16'h26c0;
assign q[5321]= 16'h2666;
assign q[5322]= 16'h2551;
assign q[5323]= 16'h238b;
assign q[5324]= 16'h2121;
assign q[5325]= 16'h1e27;
assign q[5326]= 16'h1ab5;
assign q[5327]= 16'h16e7;
assign q[5328]= 16'h12d9;
assign q[5329]= 16'heab;
assign q[5330]= 16'ha7d;
assign q[5331]= 16'h66f;
assign q[5332]= 16'h2a0;
assign q[5333]= 16'hff2d;
assign q[5334]= 16'hfc2e;
assign q[5335]= 16'hf9ba;
assign q[5336]= 16'hf7e3;
assign q[5337]= 16'hf6b8;
assign q[5338]= 16'hf641;
assign q[5339]= 16'hf684;
assign q[5340]= 16'hf77f;
assign q[5341]= 16'hf92d;
assign q[5342]= 16'hfb87;
assign q[5343]= 16'hfe7e;
assign q[5344]= 16'h201;
assign q[5345]= 16'h5ff;
assign q[5346]= 16'ha60;
assign q[5347]= 16'hf0e;
assign q[5348]= 16'h13ee;
assign q[5349]= 16'h18e9;
assign q[5350]= 16'h1de4;
assign q[5351]= 16'h22c6;
assign q[5352]= 16'h2778;
assign q[5353]= 16'h2be1;
assign q[5354]= 16'h2fec;
assign q[5355]= 16'h3387;
assign q[5356]= 16'h36a0;
assign q[5357]= 16'h3928;
assign q[5358]= 16'h3b12;
assign q[5359]= 16'h3c56;
assign q[5360]= 16'h3cec;
assign q[5361]= 16'h3ccf;
assign q[5362]= 16'h3bff;
assign q[5363]= 16'h3a7d;
assign q[5364]= 16'h384d;
assign q[5365]= 16'h3577;
assign q[5366]= 16'h3202;
assign q[5367]= 16'h2dfc;
assign q[5368]= 16'h2973;
assign q[5369]= 16'h2478;
assign q[5370]= 16'h1f1c;
assign q[5371]= 16'h1975;
assign q[5372]= 16'h1397;
assign q[5373]= 16'hd9b;
assign q[5374]= 16'h796;
assign q[5375]= 16'h1a2;
assign q[5376]= 16'hfbd7;
assign q[5377]= 16'hf64a;
assign q[5378]= 16'hf113;
assign q[5379]= 16'hec46;
assign q[5380]= 16'he7f6;
assign q[5381]= 16'he435;
assign q[5382]= 16'he110;
assign q[5383]= 16'hde94;
assign q[5384]= 16'hdcc8;
assign q[5385]= 16'hdbb1;
assign q[5386]= 16'hdb51;
assign q[5387]= 16'hdba5;
assign q[5388]= 16'hdcaa;
assign q[5389]= 16'hde55;
assign q[5390]= 16'he09c;
assign q[5391]= 16'he370;
assign q[5392]= 16'he6c0;
assign q[5393]= 16'hea7b;
assign q[5394]= 16'hee8a;
assign q[5395]= 16'hf2d9;
assign q[5396]= 16'hf751;
assign q[5397]= 16'hfbdc;
assign q[5398]= 16'h62;
assign q[5399]= 16'h4cf;
assign q[5400]= 16'h90d;
assign q[5401]= 16'hd08;
assign q[5402]= 16'h10af;
assign q[5403]= 16'h13f1;
assign q[5404]= 16'h16bf;
assign q[5405]= 16'h190f;
assign q[5406]= 16'h1ad6;
assign q[5407]= 16'h1c0d;
assign q[5408]= 16'h1cb0;
assign q[5409]= 16'h1cbc;
assign q[5410]= 16'h1c33;
assign q[5411]= 16'h1b16;
assign q[5412]= 16'h196b;
assign q[5413]= 16'h173a;
assign q[5414]= 16'h148b;
assign q[5415]= 16'h116c;
assign q[5416]= 16'hde8;
assign q[5417]= 16'ha10;
assign q[5418]= 16'h5f4;
assign q[5419]= 16'h1a6;
assign q[5420]= 16'hfd3a;
assign q[5421]= 16'hf8c1;
assign q[5422]= 16'hf44f;
assign q[5423]= 16'heffa;
assign q[5424]= 16'hebd3;
assign q[5425]= 16'he7ed;
assign q[5426]= 16'he459;
assign q[5427]= 16'he126;
assign q[5428]= 16'hde63;
assign q[5429]= 16'hdc18;
assign q[5430]= 16'hda4f;
assign q[5431]= 16'hd90c;
assign q[5432]= 16'hd851;
assign q[5433]= 16'hd81b;
assign q[5434]= 16'hd866;
assign q[5435]= 16'hd928;
assign q[5436]= 16'hda55;
assign q[5437]= 16'hdbdf;
assign q[5438]= 16'hddb3;
assign q[5439]= 16'hdfbf;
assign q[5440]= 16'he1ee;
assign q[5441]= 16'he428;
assign q[5442]= 16'he659;
assign q[5443]= 16'he86a;
assign q[5444]= 16'hea48;
assign q[5445]= 16'hebdf;
assign q[5446]= 16'hed20;
assign q[5447]= 16'hedff;
assign q[5448]= 16'hee72;
assign q[5449]= 16'hee74;
assign q[5450]= 16'hee05;
assign q[5451]= 16'hed27;
assign q[5452]= 16'hebe3;
assign q[5453]= 16'hea44;
assign q[5454]= 16'he858;
assign q[5455]= 16'he631;
assign q[5456]= 16'he3e4;
assign q[5457]= 16'he187;
assign q[5458]= 16'hdf2f;
assign q[5459]= 16'hdcf4;
assign q[5460]= 16'hdaeb;
assign q[5461]= 16'hd928;
assign q[5462]= 16'hd7bc;
assign q[5463]= 16'hd6b6;
assign q[5464]= 16'hd61f;
assign q[5465]= 16'hd5fd;
assign q[5466]= 16'hd653;
assign q[5467]= 16'hd71e;
assign q[5468]= 16'hd856;
assign q[5469]= 16'hd9f0;
assign q[5470]= 16'hdbdd;
assign q[5471]= 16'hde0b;
assign q[5472]= 16'he064;
assign q[5473]= 16'he2d1;
assign q[5474]= 16'he53d;
assign q[5475]= 16'he78f;
assign q[5476]= 16'he9b0;
assign q[5477]= 16'heb8c;
assign q[5478]= 16'hed12;
assign q[5479]= 16'hee31;
assign q[5480]= 16'heedf;
assign q[5481]= 16'hef15;
assign q[5482]= 16'heed2;
assign q[5483]= 16'hee17;
assign q[5484]= 16'hecec;
assign q[5485]= 16'heb5c;
assign q[5486]= 16'he976;
assign q[5487]= 16'he74d;
assign q[5488]= 16'he4f7;
assign q[5489]= 16'he28b;
assign q[5490]= 16'he022;
assign q[5491]= 16'hddd4;
assign q[5492]= 16'hdbbb;
assign q[5493]= 16'hd9ed;
assign q[5494]= 16'hd880;
assign q[5495]= 16'hd785;
assign q[5496]= 16'hd70e;
assign q[5497]= 16'hd723;
assign q[5498]= 16'hd7ce;
assign q[5499]= 16'hd911;
assign q[5500]= 16'hdaea;
assign q[5501]= 16'hdd56;
assign q[5502]= 16'he04a;
assign q[5503]= 16'he3ba;
assign q[5504]= 16'he797;
assign q[5505]= 16'hebcf;
assign q[5506]= 16'hf04e;
assign q[5507]= 16'hf4ff;
assign q[5508]= 16'hf9ce;
assign q[5509]= 16'hfea5;
assign q[5510]= 16'h36e;
assign q[5511]= 16'h81a;
assign q[5512]= 16'hc95;
assign q[5513]= 16'h10d1;
assign q[5514]= 16'h14c1;
assign q[5515]= 16'h185c;
assign q[5516]= 16'h1b9a;
assign q[5517]= 16'h1e77;
assign q[5518]= 16'h20f2;
assign q[5519]= 16'h230a;
assign q[5520]= 16'h24c3;
assign q[5521]= 16'h2621;
assign q[5522]= 16'h272a;
assign q[5523]= 16'h27e5;
assign q[5524]= 16'h2858;
assign q[5525]= 16'h288d;
assign q[5526]= 16'h288a;
assign q[5527]= 16'h2856;
assign q[5528]= 16'h27f8;
assign q[5529]= 16'h2775;
assign q[5530]= 16'h26d0;
assign q[5531]= 16'h260f;
assign q[5532]= 16'h2532;
assign q[5533]= 16'h243a;
assign q[5534]= 16'h2329;
assign q[5535]= 16'h21fd;
assign q[5536]= 16'h20b7;
assign q[5537]= 16'h1f55;
assign q[5538]= 16'h1dd7;
assign q[5539]= 16'h1c3d;
assign q[5540]= 16'h1a89;
assign q[5541]= 16'h18bb;
assign q[5542]= 16'h16d9;
assign q[5543]= 16'h14e6;
assign q[5544]= 16'h12e9;
assign q[5545]= 16'h10e9;
assign q[5546]= 16'hef1;
assign q[5547]= 16'hd0a;
assign q[5548]= 16'hb40;
assign q[5549]= 16'h9a0;
assign q[5550]= 16'h837;
assign q[5551]= 16'h710;
assign q[5552]= 16'h638;
assign q[5553]= 16'h5b9;
assign q[5554]= 16'h59e;
assign q[5555]= 16'h5ec;
assign q[5556]= 16'h6aa;
assign q[5557]= 16'h7d7;
assign q[5558]= 16'h974;
assign q[5559]= 16'hb7a;
assign q[5560]= 16'hde2;
assign q[5561]= 16'h109e;
assign q[5562]= 16'h13a0;
assign q[5563]= 16'h16d4;
assign q[5564]= 16'h1a25;
assign q[5565]= 16'h1d7c;
assign q[5566]= 16'h20be;
assign q[5567]= 16'h23d2;
assign q[5568]= 16'h269d;
assign q[5569]= 16'h2904;
assign q[5570]= 16'h2af0;
assign q[5571]= 16'h2c4a;
assign q[5572]= 16'h2d00;
assign q[5573]= 16'h2d01;
assign q[5574]= 16'h2c43;
assign q[5575]= 16'h2ac0;
assign q[5576]= 16'h2878;
assign q[5577]= 16'h256f;
assign q[5578]= 16'h21ae;
assign q[5579]= 16'h1d47;
assign q[5580]= 16'h184c;
assign q[5581]= 16'h12d7;
assign q[5582]= 16'hd04;
assign q[5583]= 16'h6f2;
assign q[5584]= 16'hc3;
assign q[5585]= 16'hfa9a;
assign q[5586]= 16'hf498;
assign q[5587]= 16'heede;
assign q[5588]= 16'he98b;
assign q[5589]= 16'he4bc;
assign q[5590]= 16'he087;
assign q[5591]= 16'hdd01;
assign q[5592]= 16'hda35;
assign q[5593]= 16'hd82d;
assign q[5594]= 16'hd6ea;
assign q[5595]= 16'hd667;
assign q[5596]= 16'hd69a;
assign q[5597]= 16'hd774;
assign q[5598]= 16'hd8e0;
assign q[5599]= 16'hdac5;
assign q[5600]= 16'hdd09;
assign q[5601]= 16'hdf8c;
assign q[5602]= 16'he230;
assign q[5603]= 16'he4d6;
assign q[5604]= 16'he75e;
assign q[5605]= 16'he9af;
assign q[5606]= 16'hebad;
assign q[5607]= 16'hed46;
assign q[5608]= 16'hee68;
assign q[5609]= 16'hef07;
assign q[5610]= 16'hef20;
assign q[5611]= 16'heeb1;
assign q[5612]= 16'hedc0;
assign q[5613]= 16'hec58;
assign q[5614]= 16'hea89;
assign q[5615]= 16'he866;
assign q[5616]= 16'he608;
assign q[5617]= 16'he387;
assign q[5618]= 16'he100;
assign q[5619]= 16'hde8e;
assign q[5620]= 16'hdc4e;
assign q[5621]= 16'hda59;
assign q[5622]= 16'hd8c7;
assign q[5623]= 16'hd7ae;
assign q[5624]= 16'hd71e;
assign q[5625]= 16'hd724;
assign q[5626]= 16'hd7c9;
assign q[5627]= 16'hd90e;
assign q[5628]= 16'hdaf3;
assign q[5629]= 16'hdd70;
assign q[5630]= 16'he07b;
assign q[5631]= 16'he404;
assign q[5632]= 16'he7f8;
assign q[5633]= 16'hec41;
assign q[5634]= 16'hf0c9;
assign q[5635]= 16'hf576;
assign q[5636]= 16'hfa2e;
assign q[5637]= 16'hfed9;
assign q[5638]= 16'h35c;
assign q[5639]= 16'h7a4;
assign q[5640]= 16'hb9b;
assign q[5641]= 16'hf30;
assign q[5642]= 16'h1253;
assign q[5643]= 16'h14f8;
assign q[5644]= 16'h1719;
assign q[5645]= 16'h18b1;
assign q[5646]= 16'h19bd;
assign q[5647]= 16'h1a3f;
assign q[5648]= 16'h1a3c;
assign q[5649]= 16'h19b9;
assign q[5650]= 16'h18c0;
assign q[5651]= 16'h1759;
assign q[5652]= 16'h1591;
assign q[5653]= 16'h1371;
assign q[5654]= 16'h1106;
assign q[5655]= 16'he5c;
assign q[5656]= 16'hb7d;
assign q[5657]= 16'h874;
assign q[5658]= 16'h54a;
assign q[5659]= 16'h209;
assign q[5660]= 16'hfeb8;
assign q[5661]= 16'hfb5d;
assign q[5662]= 16'hf800;
assign q[5663]= 16'hf4a6;
assign q[5664]= 16'hf154;
assign q[5665]= 16'hee10;
assign q[5666]= 16'heae0;
assign q[5667]= 16'he7c8;
assign q[5668]= 16'he4cf;
assign q[5669]= 16'he1fb;
assign q[5670]= 16'hdf54;
assign q[5671]= 16'hdce2;
assign q[5672]= 16'hdaac;
assign q[5673]= 16'hd8bc;
assign q[5674]= 16'hd71b;
assign q[5675]= 16'hd5d3;
assign q[5676]= 16'hd4ed;
assign q[5677]= 16'hd473;
assign q[5678]= 16'hd46c;
assign q[5679]= 16'hd4e0;
assign q[5680]= 16'hd5d5;
assign q[5681]= 16'hd74d;
assign q[5682]= 16'hd94c;
assign q[5683]= 16'hdbd1;
assign q[5684]= 16'hded8;
assign q[5685]= 16'he25b;
assign q[5686]= 16'he652;
assign q[5687]= 16'heab0;
assign q[5688]= 16'hef66;
assign q[5689]= 16'hf465;
assign q[5690]= 16'hf997;
assign q[5691]= 16'hfee7;
assign q[5692]= 16'h43e;
assign q[5693]= 16'h984;
assign q[5694]= 16'hea1;
assign q[5695]= 16'h137b;
assign q[5696]= 16'h17fb;
assign q[5697]= 16'h1c0a;
assign q[5698]= 16'h1f93;
assign q[5699]= 16'h2286;
assign q[5700]= 16'h24d3;
assign q[5701]= 16'h2670;
assign q[5702]= 16'h2755;
assign q[5703]= 16'h277f;
assign q[5704]= 16'h26f1;
assign q[5705]= 16'h25b1;
assign q[5706]= 16'h23c9;
assign q[5707]= 16'h214a;
assign q[5708]= 16'h1e45;
assign q[5709]= 16'h1ad2;
assign q[5710]= 16'h170a;
assign q[5711]= 16'h1309;
assign q[5712]= 16'heed;
assign q[5713]= 16'had3;
assign q[5714]= 16'h6da;
assign q[5715]= 16'h320;
assign q[5716]= 16'hffc0;
assign q[5717]= 16'hfcd3;
assign q[5718]= 16'hfa6e;
assign q[5719]= 16'hf8a4;
assign q[5720]= 16'hf784;
assign q[5721]= 16'hf715;
assign q[5722]= 16'hf75d;
assign q[5723]= 16'hf85a;
assign q[5724]= 16'hfa07;
assign q[5725]= 16'hfc59;
assign q[5726]= 16'hff40;
assign q[5727]= 16'h2a9;
assign q[5728]= 16'h681;
assign q[5729]= 16'haac;
assign q[5730]= 16'hf10;
assign q[5731]= 16'h1392;
assign q[5732]= 16'h1817;
assign q[5733]= 16'h1c83;
assign q[5734]= 16'h20bd;
assign q[5735]= 16'h24af;
assign q[5736]= 16'h2845;
assign q[5737]= 16'h2b6e;
assign q[5738]= 16'h2e1f;
assign q[5739]= 16'h3050;
assign q[5740]= 16'h31fc;
assign q[5741]= 16'h3326;
assign q[5742]= 16'h33d3;
assign q[5743]= 16'h340a;
assign q[5744]= 16'h33d8;
assign q[5745]= 16'h334c;
assign q[5746]= 16'h3278;
assign q[5747]= 16'h316d;
assign q[5748]= 16'h303e;
assign q[5749]= 16'h2eff;
assign q[5750]= 16'h2dc1;
assign q[5751]= 16'h2c94;
assign q[5752]= 16'h2b87;
assign q[5753]= 16'h2aa5;
assign q[5754]= 16'h29f7;
assign q[5755]= 16'h2981;
assign q[5756]= 16'h2946;
assign q[5757]= 16'h2943;
assign q[5758]= 16'h2973;
assign q[5759]= 16'h29d1;
assign q[5760]= 16'h2a50;
assign q[5761]= 16'h2ae5;
assign q[5762]= 16'h2b83;
assign q[5763]= 16'h2c1c;
assign q[5764]= 16'h2ca2;
assign q[5765]= 16'h2d07;
assign q[5766]= 16'h2d3e;
assign q[5767]= 16'h2d3d;
assign q[5768]= 16'h2cfb;
assign q[5769]= 16'h2c72;
assign q[5770]= 16'h2b9f;
assign q[5771]= 16'h2a80;
assign q[5772]= 16'h2918;
assign q[5773]= 16'h276b;
assign q[5774]= 16'h257f;
assign q[5775]= 16'h235f;
assign q[5776]= 16'h2113;
assign q[5777]= 16'h1ea8;
assign q[5778]= 16'h1c29;
assign q[5779]= 16'h19a3;
assign q[5780]= 16'h1720;
assign q[5781]= 16'h14ab;
assign q[5782]= 16'h124c;
assign q[5783]= 16'h100a;
assign q[5784]= 16'hdeb;
assign q[5785]= 16'hbf0;
assign q[5786]= 16'ha1b;
assign q[5787]= 16'h869;
assign q[5788]= 16'h6d7;
assign q[5789]= 16'h55f;
assign q[5790]= 16'h3fb;
assign q[5791]= 16'h2a3;
assign q[5792]= 16'h150;
assign q[5793]= 16'hfffa;
assign q[5794]= 16'hfe99;
assign q[5795]= 16'hfd28;
assign q[5796]= 16'hfba3;
assign q[5797]= 16'hfa07;
assign q[5798]= 16'hf854;
assign q[5799]= 16'hf68d;
assign q[5800]= 16'hf4b6;
assign q[5801]= 16'hf2d7;
assign q[5802]= 16'hf0f9;
assign q[5803]= 16'hef27;
assign q[5804]= 16'hed6f;
assign q[5805]= 16'hebde;
assign q[5806]= 16'hea83;
assign q[5807]= 16'he96d;
assign q[5808]= 16'he8a9;
assign q[5809]= 16'he845;
assign q[5810]= 16'he84c;
assign q[5811]= 16'he8c7;
assign q[5812]= 16'he9bc;
assign q[5813]= 16'heb2d;
assign q[5814]= 16'hed1c;
assign q[5815]= 16'hef84;
assign q[5816]= 16'hf25f;
assign q[5817]= 16'hf5a1;
assign q[5818]= 16'hf93f;
assign q[5819]= 16'hfd26;
assign q[5820]= 16'h144;
assign q[5821]= 16'h586;
assign q[5822]= 16'h9d6;
assign q[5823]= 16'he1b;
assign q[5824]= 16'h1240;
assign q[5825]= 16'h162f;
assign q[5826]= 16'h19d2;
assign q[5827]= 16'h1d15;
assign q[5828]= 16'h1fe7;
assign q[5829]= 16'h223a;
assign q[5830]= 16'h2401;
assign q[5831]= 16'h2534;
assign q[5832]= 16'h25cd;
assign q[5833]= 16'h25ca;
assign q[5834]= 16'h252c;
assign q[5835]= 16'h23f8;
assign q[5836]= 16'h2236;
assign q[5837]= 16'h1fef;
assign q[5838]= 16'h1d30;
assign q[5839]= 16'h1a09;
assign q[5840]= 16'h1688;
assign q[5841]= 16'h12c1;
assign q[5842]= 16'hec6;
assign q[5843]= 16'haa9;
assign q[5844]= 16'h67e;
assign q[5845]= 16'h257;
assign q[5846]= 16'hfe48;
assign q[5847]= 16'hfa5f;
assign q[5848]= 16'hf6ad;
assign q[5849]= 16'hf342;
assign q[5850]= 16'hf029;
assign q[5851]= 16'hed6e;
assign q[5852]= 16'heb1a;
assign q[5853]= 16'he934;
assign q[5854]= 16'he7c2;
assign q[5855]= 16'he6c8;
assign q[5856]= 16'he645;
assign q[5857]= 16'he639;
assign q[5858]= 16'he6a2;
assign q[5859]= 16'he77a;
assign q[5860]= 16'he8ba;
assign q[5861]= 16'hea5b;
assign q[5862]= 16'hec51;
assign q[5863]= 16'hee92;
assign q[5864]= 16'hf110;
assign q[5865]= 16'hf3bd;
assign q[5866]= 16'hf68a;
assign q[5867]= 16'hf967;
assign q[5868]= 16'hfc45;
assign q[5869]= 16'hff13;
assign q[5870]= 16'h1c0;
assign q[5871]= 16'h440;
assign q[5872]= 16'h684;
assign q[5873]= 16'h87f;
assign q[5874]= 16'ha26;
assign q[5875]= 16'hb70;
assign q[5876]= 16'hc57;
assign q[5877]= 16'hcd6;
assign q[5878]= 16'hced;
assign q[5879]= 16'hc9c;
assign q[5880]= 16'hbe7;
assign q[5881]= 16'had5;
assign q[5882]= 16'h971;
assign q[5883]= 16'h7c4;
assign q[5884]= 16'h5df;
assign q[5885]= 16'h3cf;
assign q[5886]= 16'h1a7;
assign q[5887]= 16'hff7a;
assign q[5888]= 16'hfd58;
assign q[5889]= 16'hfb55;
assign q[5890]= 16'hf983;
assign q[5891]= 16'hf7f3;
assign q[5892]= 16'hf6b4;
assign q[5893]= 16'hf5d4;
assign q[5894]= 16'hf55e;
assign q[5895]= 16'hf55b;
assign q[5896]= 16'hf5d1;
assign q[5897]= 16'hf6c2;
assign q[5898]= 16'hf82d;
assign q[5899]= 16'hfa10;
assign q[5900]= 16'hfc64;
assign q[5901]= 16'hff21;
assign q[5902]= 16'h238;
assign q[5903]= 16'h5a0;
assign q[5904]= 16'h947;
assign q[5905]= 16'hd1d;
assign q[5906]= 16'h1110;
assign q[5907]= 16'h150e;
assign q[5908]= 16'h1905;
assign q[5909]= 16'h1ce5;
assign q[5910]= 16'h209d;
assign q[5911]= 16'h241e;
assign q[5912]= 16'h275a;
assign q[5913]= 16'h2a47;
assign q[5914]= 16'h2cdb;
assign q[5915]= 16'h2f0f;
assign q[5916]= 16'h30df;
assign q[5917]= 16'h3249;
assign q[5918]= 16'h334d;
assign q[5919]= 16'h33ed;
assign q[5920]= 16'h342f;
assign q[5921]= 16'h341a;
assign q[5922]= 16'h33b4;
assign q[5923]= 16'h3309;
assign q[5924]= 16'h3222;
assign q[5925]= 16'h310d;
assign q[5926]= 16'h2fd4;
assign q[5927]= 16'h2e86;
assign q[5928]= 16'h2d2d;
assign q[5929]= 16'h2bd7;
assign q[5930]= 16'h2a8f;
assign q[5931]= 16'h2960;
assign q[5932]= 16'h2854;
assign q[5933]= 16'h2773;
assign q[5934]= 16'h26c5;
assign q[5935]= 16'h264e;
assign q[5936]= 16'h2614;
assign q[5937]= 16'h2619;
assign q[5938]= 16'h265b;
assign q[5939]= 16'h26db;
assign q[5940]= 16'h2795;
assign q[5941]= 16'h2883;
assign q[5942]= 16'h299e;
assign q[5943]= 16'h2adf;
assign q[5944]= 16'h2c3b;
assign q[5945]= 16'h2da6;
assign q[5946]= 16'h2f15;
assign q[5947]= 16'h307a;
assign q[5948]= 16'h31c8;
assign q[5949]= 16'h32ef;
assign q[5950]= 16'h33e3;
assign q[5951]= 16'h3494;
assign q[5952]= 16'h34f7;
assign q[5953]= 16'h3500;
assign q[5954]= 16'h34a2;
assign q[5955]= 16'h33d7;
assign q[5956]= 16'h3295;
assign q[5957]= 16'h30d9;
assign q[5958]= 16'h2ea0;
assign q[5959]= 16'h2be9;
assign q[5960]= 16'h28b7;
assign q[5961]= 16'h250f;
assign q[5962]= 16'h20f8;
assign q[5963]= 16'h1c7d;
assign q[5964]= 16'h17aa;
assign q[5965]= 16'h128d;
assign q[5966]= 16'hd37;
assign q[5967]= 16'h7b9;
assign q[5968]= 16'h227;
assign q[5969]= 16'hfc95;
assign q[5970]= 16'hf716;
assign q[5971]= 16'hf1be;
assign q[5972]= 16'heca2;
assign q[5973]= 16'he7d3;
assign q[5974]= 16'he365;
assign q[5975]= 16'hdf66;
assign q[5976]= 16'hdbe6;
assign q[5977]= 16'hd8ef;
assign q[5978]= 16'hd68c;
assign q[5979]= 16'hd4c4;
assign q[5980]= 16'hd39c;
assign q[5981]= 16'hd314;
assign q[5982]= 16'hd32c;
assign q[5983]= 16'hd3e0;
assign q[5984]= 16'hd52b;
assign q[5985]= 16'hd702;
assign q[5986]= 16'hd95c;
assign q[5987]= 16'hdc2b;
assign q[5988]= 16'hdf60;
assign q[5989]= 16'he2eb;
assign q[5990]= 16'he6ba;
assign q[5991]= 16'heaba;
assign q[5992]= 16'heed7;
assign q[5993]= 16'hf2ff;
assign q[5994]= 16'hf71d;
assign q[5995]= 16'hfb1d;
assign q[5996]= 16'hfeed;
assign q[5997]= 16'h27a;
assign q[5998]= 16'h5b4;
assign q[5999]= 16'h88c;
assign q[6000]= 16'haf4;
assign q[6001]= 16'hce0;
assign q[6002]= 16'he48;
assign q[6003]= 16'hf24;
assign q[6004]= 16'hf71;
assign q[6005]= 16'hf2d;
assign q[6006]= 16'he5a;
assign q[6007]= 16'hcfc;
assign q[6008]= 16'hb1b;
assign q[6009]= 16'h8bf;
assign q[6010]= 16'h5f5;
assign q[6011]= 16'h2cd;
assign q[6012]= 16'hff57;
assign q[6013]= 16'hfba3;
assign q[6014]= 16'hf7c8;
assign q[6015]= 16'hf3d8;
assign q[6016]= 16'hefea;
assign q[6017]= 16'hec10;
assign q[6018]= 16'he861;
assign q[6019]= 16'he4ef;
assign q[6020]= 16'he1ca;
assign q[6021]= 16'hdf03;
assign q[6022]= 16'hdca6;
assign q[6023]= 16'hdabd;
assign q[6024]= 16'hd950;
assign q[6025]= 16'hd861;
assign q[6026]= 16'hd7f2;
assign q[6027]= 16'hd7fe;
assign q[6028]= 16'hd880;
assign q[6029]= 16'hd96e;
assign q[6030]= 16'hdabc;
assign q[6031]= 16'hdc5b;
assign q[6032]= 16'hde3a;
assign q[6033]= 16'he047;
assign q[6034]= 16'he270;
assign q[6035]= 16'he49f;
assign q[6036]= 16'he6c2;
assign q[6037]= 16'he8c7;
assign q[6038]= 16'hea9b;
assign q[6039]= 16'hec2e;
assign q[6040]= 16'hed74;
assign q[6041]= 16'hee62;
assign q[6042]= 16'heeee;
assign q[6043]= 16'hef14;
assign q[6044]= 16'heed1;
assign q[6045]= 16'hee26;
assign q[6046]= 16'hed18;
assign q[6047]= 16'hebab;
assign q[6048]= 16'he9e9;
assign q[6049]= 16'he7dd;
assign q[6050]= 16'he594;
assign q[6051]= 16'he31c;
assign q[6052]= 16'he084;
assign q[6053]= 16'hdddc;
assign q[6054]= 16'hdb32;
assign q[6055]= 16'hd898;
assign q[6056]= 16'hd61a;
assign q[6057]= 16'hd3c6;
assign q[6058]= 16'hd1a9;
assign q[6059]= 16'hcfce;
assign q[6060]= 16'hce3c;
assign q[6061]= 16'hccfb;
assign q[6062]= 16'hcc10;
assign q[6063]= 16'hcb7f;
assign q[6064]= 16'hcb47;
assign q[6065]= 16'hcb6a;
assign q[6066]= 16'hcbe4;
assign q[6067]= 16'hccb1;
assign q[6068]= 16'hcdcd;
assign q[6069]= 16'hcf31;
assign q[6070]= 16'hd0d4;
assign q[6071]= 16'hd2af;
assign q[6072]= 16'hd4b8;
assign q[6073]= 16'hd6e5;
assign q[6074]= 16'hd92c;
assign q[6075]= 16'hdb82;
assign q[6076]= 16'hdddc;
assign q[6077]= 16'he02f;
assign q[6078]= 16'he270;
assign q[6079]= 16'he496;
assign q[6080]= 16'he696;
assign q[6081]= 16'he867;
assign q[6082]= 16'hea01;
assign q[6083]= 16'heb5c;
assign q[6084]= 16'hec73;
assign q[6085]= 16'hed3f;
assign q[6086]= 16'hedbd;
assign q[6087]= 16'hedeb;
assign q[6088]= 16'hedca;
assign q[6089]= 16'hed5a;
assign q[6090]= 16'hec9e;
assign q[6091]= 16'heb9b;
assign q[6092]= 16'hea59;
assign q[6093]= 16'he8de;
assign q[6094]= 16'he736;
assign q[6095]= 16'he56b;
assign q[6096]= 16'he388;
assign q[6097]= 16'he19c;
assign q[6098]= 16'hdfb3;
assign q[6099]= 16'hdddb;
assign q[6100]= 16'hdc21;
assign q[6101]= 16'hda91;
assign q[6102]= 16'hd938;
assign q[6103]= 16'hd81f;
assign q[6104]= 16'hd750;
assign q[6105]= 16'hd6d1;
assign q[6106]= 16'hd6a7;
assign q[6107]= 16'hd6d5;
assign q[6108]= 16'hd75c;
assign q[6109]= 16'hd839;
assign q[6110]= 16'hd968;
assign q[6111]= 16'hdae4;
assign q[6112]= 16'hdca4;
assign q[6113]= 16'hde9e;
assign q[6114]= 16'he0c8;
assign q[6115]= 16'he316;
assign q[6116]= 16'he57a;
assign q[6117]= 16'he7e7;
assign q[6118]= 16'hea51;
assign q[6119]= 16'hecaa;
assign q[6120]= 16'heee6;
assign q[6121]= 16'hf0fb;
assign q[6122]= 16'hf2de;
assign q[6123]= 16'hf486;
assign q[6124]= 16'hf5ed;
assign q[6125]= 16'hf70c;
assign q[6126]= 16'hf7df;
assign q[6127]= 16'hf864;
assign q[6128]= 16'hf89a;
assign q[6129]= 16'hf882;
assign q[6130]= 16'hf81c;
assign q[6131]= 16'hf76c;
assign q[6132]= 16'hf676;
assign q[6133]= 16'hf53f;
assign q[6134]= 16'hf3cd;
assign q[6135]= 16'hf226;
assign q[6136]= 16'hf052;
assign q[6137]= 16'hee59;
assign q[6138]= 16'hec42;
assign q[6139]= 16'hea16;
assign q[6140]= 16'he7df;
assign q[6141]= 16'he5a6;
assign q[6142]= 16'he373;
assign q[6143]= 16'he151;
assign q[6144]= 16'hdf48;
assign q[6145]= 16'hdd63;
assign q[6146]= 16'hdbaa;
assign q[6147]= 16'hda26;
assign q[6148]= 16'hd8df;
assign q[6149]= 16'hd7dd;
assign q[6150]= 16'hd725;
assign q[6151]= 16'hd6bb;
assign q[6152]= 16'hd6a4;
assign q[6153]= 16'hd6e1;
assign q[6154]= 16'hd771;
assign q[6155]= 16'hd853;
assign q[6156]= 16'hd981;
assign q[6157]= 16'hdaf4;
assign q[6158]= 16'hdca5;
assign q[6159]= 16'hde8a;
assign q[6160]= 16'he095;
assign q[6161]= 16'he2b9;
assign q[6162]= 16'he4e9;
assign q[6163]= 16'he716;
assign q[6164]= 16'he931;
assign q[6165]= 16'heb2c;
assign q[6166]= 16'hecfa;
assign q[6167]= 16'hee91;
assign q[6168]= 16'hefe7;
assign q[6169]= 16'hf0f6;
assign q[6170]= 16'hf1bb;
assign q[6171]= 16'hf235;
assign q[6172]= 16'hf268;
assign q[6173]= 16'hf259;
assign q[6174]= 16'hf213;
assign q[6175]= 16'hf1a1;
assign q[6176]= 16'hf112;
assign q[6177]= 16'hf077;
assign q[6178]= 16'hefe1;
assign q[6179]= 16'hef62;
assign q[6180]= 16'hef0c;
assign q[6181]= 16'heeef;
assign q[6182]= 16'hef19;
assign q[6183]= 16'hef95;
assign q[6184]= 16'hf06d;
assign q[6185]= 16'hf1a3;
assign q[6186]= 16'hf338;
assign q[6187]= 16'hf526;
assign q[6188]= 16'hf766;
assign q[6189]= 16'hf9e8;
assign q[6190]= 16'hfc9c;
assign q[6191]= 16'hff6d;
assign q[6192]= 16'h243;
assign q[6193]= 16'h505;
assign q[6194]= 16'h79b;
assign q[6195]= 16'h9ea;
assign q[6196]= 16'hbdb;
assign q[6197]= 16'hd5a;
assign q[6198]= 16'he54;
assign q[6199]= 16'hebe;
assign q[6200]= 16'he91;
assign q[6201]= 16'hdcb;
assign q[6202]= 16'hc70;
assign q[6203]= 16'ha8e;
assign q[6204]= 16'h834;
assign q[6205]= 16'h57a;
assign q[6206]= 16'h27c;
assign q[6207]= 16'hff5a;
assign q[6208]= 16'hfc35;
assign q[6209]= 16'hf932;
assign q[6210]= 16'hf676;
assign q[6211]= 16'hf422;
assign q[6212]= 16'hf256;
assign q[6213]= 16'hf12e;
assign q[6214]= 16'hf0c0;
assign q[6215]= 16'hf11b;
assign q[6216]= 16'hf247;
assign q[6217]= 16'hf443;
assign q[6218]= 16'hf707;
assign q[6219]= 16'hfa84;
assign q[6220]= 16'hfea0;
assign q[6221]= 16'h33b;
assign q[6222]= 16'h832;
assign q[6223]= 16'hd59;
assign q[6224]= 16'h1284;
assign q[6225]= 16'h1783;
assign q[6226]= 16'h1c27;
assign q[6227]= 16'h2043;
assign q[6228]= 16'h23ad;
assign q[6229]= 16'h2642;
assign q[6230]= 16'h27e4;
assign q[6231]= 16'h287c;
assign q[6232]= 16'h27fe;
assign q[6233]= 16'h2666;
assign q[6234]= 16'h23ba;
assign q[6235]= 16'h2009;
assign q[6236]= 16'h1b6c;
assign q[6237]= 16'h1603;
assign q[6238]= 16'hff7;
assign q[6239]= 16'h974;
assign q[6240]= 16'h2ac;
assign q[6241]= 16'hfbd5;
assign q[6242]= 16'hf520;
assign q[6243]= 16'heec1;
assign q[6244]= 16'he8e9;
assign q[6245]= 16'he3c2;
assign q[6246]= 16'hdf70;
assign q[6247]= 16'hdc12;
assign q[6248]= 16'hd9bb;
assign q[6249]= 16'hd877;
assign q[6250]= 16'hd847;
assign q[6251]= 16'hd924;
assign q[6252]= 16'hdaff;
assign q[6253]= 16'hddbd;
assign q[6254]= 16'he141;
assign q[6255]= 16'he563;
assign q[6256]= 16'he9fa;
assign q[6257]= 16'heedb;
assign q[6258]= 16'hf3d6;
assign q[6259]= 16'hf8bf;
assign q[6260]= 16'hfd6b;
assign q[6261]= 16'h1b2;
assign q[6262]= 16'h575;
assign q[6263]= 16'h896;
assign q[6264]= 16'hb02;
assign q[6265]= 16'hcac;
assign q[6266]= 16'hd8e;
assign q[6267]= 16'hdac;
assign q[6268]= 16'hd10;
assign q[6269]= 16'hbcc;
assign q[6270]= 16'h9f7;
assign q[6271]= 16'h7ae;
assign q[6272]= 16'h511;
assign q[6273]= 16'h242;
assign q[6274]= 16'hff68;
assign q[6275]= 16'hfca2;
assign q[6276]= 16'hfa16;
assign q[6277]= 16'hf7e2;
assign q[6278]= 16'hf621;
assign q[6279]= 16'hf4eb;
assign q[6280]= 16'hf452;
assign q[6281]= 16'hf461;
assign q[6282]= 16'hf51d;
assign q[6283]= 16'hf688;
assign q[6284]= 16'hf89b;
assign q[6285]= 16'hfb4b;
assign q[6286]= 16'hfe88;
assign q[6287]= 16'h23d;
assign q[6288]= 16'h655;
assign q[6289]= 16'hab5;
assign q[6290]= 16'hf44;
assign q[6291]= 16'h13e6;
assign q[6292]= 16'h1881;
assign q[6293]= 16'h1cfc;
assign q[6294]= 16'h2140;
assign q[6295]= 16'h2539;
assign q[6296]= 16'h28d6;
assign q[6297]= 16'h2c09;
assign q[6298]= 16'h2ec8;
assign q[6299]= 16'h310d;
assign q[6300]= 16'h32d6;
assign q[6301]= 16'h3422;
assign q[6302]= 16'h34f5;
assign q[6303]= 16'h3555;
assign q[6304]= 16'h354b;
assign q[6305]= 16'h34e1;
assign q[6306]= 16'h3421;
assign q[6307]= 16'h3317;
assign q[6308]= 16'h31cf;
assign q[6309]= 16'h3055;
assign q[6310]= 16'h2eb4;
assign q[6311]= 16'h2cf7;
assign q[6312]= 16'h2b26;
assign q[6313]= 16'h294a;
assign q[6314]= 16'h276a;
assign q[6315]= 16'h258b;
assign q[6316]= 16'h23b1;
assign q[6317]= 16'h21e0;
assign q[6318]= 16'h2018;
assign q[6319]= 16'h1e5c;
assign q[6320]= 16'h1caa;
assign q[6321]= 16'h1b04;
assign q[6322]= 16'h1967;
assign q[6323]= 16'h17d2;
assign q[6324]= 16'h1644;
assign q[6325]= 16'h14bb;
assign q[6326]= 16'h1334;
assign q[6327]= 16'h11ae;
assign q[6328]= 16'h1028;
assign q[6329]= 16'he9e;
assign q[6330]= 16'hd0f;
assign q[6331]= 16'hb79;
assign q[6332]= 16'h9da;
assign q[6333]= 16'h830;
assign q[6334]= 16'h67b;
assign q[6335]= 16'h4b7;
assign q[6336]= 16'h2e3;
assign q[6337]= 16'hff;
assign q[6338]= 16'hff09;
assign q[6339]= 16'hfd00;
assign q[6340]= 16'hfae3;
assign q[6341]= 16'hf8b4;
assign q[6342]= 16'hf673;
assign q[6343]= 16'hf422;
assign q[6344]= 16'hf1c3;
assign q[6345]= 16'hef5a;
assign q[6346]= 16'hecea;
assign q[6347]= 16'hea7a;
assign q[6348]= 16'he80f;
assign q[6349]= 16'he5b0;
assign q[6350]= 16'he364;
assign q[6351]= 16'he135;
assign q[6352]= 16'hdf2a;
assign q[6353]= 16'hdd4c;
assign q[6354]= 16'hdba5;
assign q[6355]= 16'hda3e;
assign q[6356]= 16'hd91f;
assign q[6357]= 16'hd851;
assign q[6358]= 16'hd7da;
assign q[6359]= 16'hd7c2;
assign q[6360]= 16'hd80d;
assign q[6361]= 16'hd8bf;
assign q[6362]= 16'hd9da;
assign q[6363]= 16'hdb60;
assign q[6364]= 16'hdd4f;
assign q[6365]= 16'hdfa5;
assign q[6366]= 16'he25e;
assign q[6367]= 16'he574;
assign q[6368]= 16'he8df;
assign q[6369]= 16'hec96;
assign q[6370]= 16'hf090;
assign q[6371]= 16'hf4c1;
assign q[6372]= 16'hf91d;
assign q[6373]= 16'hfd96;
assign q[6374]= 16'h21e;
assign q[6375]= 16'h6a9;
assign q[6376]= 16'hb27;
assign q[6377]= 16'hf8a;
assign q[6378]= 16'h13c4;
assign q[6379]= 16'h17c8;
assign q[6380]= 16'h1b89;
assign q[6381]= 16'h1efb;
assign q[6382]= 16'h2214;
assign q[6383]= 16'h24c9;
assign q[6384]= 16'h2712;
assign q[6385]= 16'h28e9;
assign q[6386]= 16'h2a49;
assign q[6387]= 16'h2b2d;
assign q[6388]= 16'h2b95;
assign q[6389]= 16'h2b81;
assign q[6390]= 16'h2af1;
assign q[6391]= 16'h29eb;
assign q[6392]= 16'h2873;
assign q[6393]= 16'h268f;
assign q[6394]= 16'h2449;
assign q[6395]= 16'h21aa;
assign q[6396]= 16'h1ebe;
assign q[6397]= 16'h1b8f;
assign q[6398]= 16'h182a;
assign q[6399]= 16'h149e;
assign q[6400]= 16'h10f7;
assign q[6401]= 16'hd43;
assign q[6402]= 16'h990;
assign q[6403]= 16'h5eb;
assign q[6404]= 16'h260;
assign q[6405]= 16'hfefc;
assign q[6406]= 16'hfbc8;
assign q[6407]= 16'hf8ce;
assign q[6408]= 16'hf615;
assign q[6409]= 16'hf3a4;
assign q[6410]= 16'hf181;
assign q[6411]= 16'hefaf;
assign q[6412]= 16'hee2e;
assign q[6413]= 16'hed00;
assign q[6414]= 16'hec23;
assign q[6415]= 16'heb94;
assign q[6416]= 16'heb4f;
assign q[6417]= 16'heb4e;
assign q[6418]= 16'heb8c;
assign q[6419]= 16'hec00;
assign q[6420]= 16'heca4;
assign q[6421]= 16'hed6e;
assign q[6422]= 16'hee55;
assign q[6423]= 16'hef51;
assign q[6424]= 16'hf058;
assign q[6425]= 16'hf161;
assign q[6426]= 16'hf263;
assign q[6427]= 16'hf357;
assign q[6428]= 16'hf434;
assign q[6429]= 16'hf4f3;
assign q[6430]= 16'hf58e;
assign q[6431]= 16'hf5fe;
assign q[6432]= 16'hf63f;
assign q[6433]= 16'hf64d;
assign q[6434]= 16'hf626;
assign q[6435]= 16'hf5c6;
assign q[6436]= 16'hf52e;
assign q[6437]= 16'hf45e;
assign q[6438]= 16'hf356;
assign q[6439]= 16'hf21a;
assign q[6440]= 16'hf0ae;
assign q[6441]= 16'hef15;
assign q[6442]= 16'hed55;
assign q[6443]= 16'heb75;
assign q[6444]= 16'he97c;
assign q[6445]= 16'he772;
assign q[6446]= 16'he55f;
assign q[6447]= 16'he34b;
assign q[6448]= 16'he13f;
assign q[6449]= 16'hdf43;
assign q[6450]= 16'hdd5f;
assign q[6451]= 16'hdb9b;
assign q[6452]= 16'hd9fd;
assign q[6453]= 16'hd88b;
assign q[6454]= 16'hd748;
assign q[6455]= 16'hd638;
assign q[6456]= 16'hd55b;
assign q[6457]= 16'hd4b1;
assign q[6458]= 16'hd439;
assign q[6459]= 16'hd3ee;
assign q[6460]= 16'hd3cc;
assign q[6461]= 16'hd3cc;
assign q[6462]= 16'hd3e7;
assign q[6463]= 16'hd415;
assign q[6464]= 16'hd44d;
assign q[6465]= 16'hd487;
assign q[6466]= 16'hd4ba;
assign q[6467]= 16'hd4dd;
assign q[6468]= 16'hd4ea;
assign q[6469]= 16'hd4db;
assign q[6470]= 16'hd4ac;
assign q[6471]= 16'hd45b;
assign q[6472]= 16'hd3e8;
assign q[6473]= 16'hd355;
assign q[6474]= 16'hd2a7;
assign q[6475]= 16'hd1e4;
assign q[6476]= 16'hd116;
assign q[6477]= 16'hd047;
assign q[6478]= 16'hcf84;
assign q[6479]= 16'hcedb;
assign q[6480]= 16'hce5a;
assign q[6481]= 16'hce10;
assign q[6482]= 16'hce0d;
assign q[6483]= 16'hce5f;
assign q[6484]= 16'hcf12;
assign q[6485]= 16'hd033;
assign q[6486]= 16'hd1ca;
assign q[6487]= 16'hd3de;
assign q[6488]= 16'hd673;
assign q[6489]= 16'hd98b;
assign q[6490]= 16'hdd22;
assign q[6491]= 16'he133;
assign q[6492]= 16'he5b5;
assign q[6493]= 16'hea9d;
assign q[6494]= 16'hefdb;
assign q[6495]= 16'hf560;
assign q[6496]= 16'hfb17;
assign q[6497]= 16'hed;
assign q[6498]= 16'h6cd;
assign q[6499]= 16'hca1;
assign q[6500]= 16'h1254;
assign q[6501]= 16'h17d0;
assign q[6502]= 16'h1d04;
assign q[6503]= 16'h21dc;
assign q[6504]= 16'h264a;
assign q[6505]= 16'h2a41;
assign q[6506]= 16'h2db6;
assign q[6507]= 16'h30a2;
assign q[6508]= 16'h3301;
assign q[6509]= 16'h34d1;
assign q[6510]= 16'h3614;
assign q[6511]= 16'h36cc;
assign q[6512]= 16'h3702;
assign q[6513]= 16'h36bd;
assign q[6514]= 16'h3608;
assign q[6515]= 16'h34ee;
assign q[6516]= 16'h337d;
assign q[6517]= 16'h31c1;
assign q[6518]= 16'h2fc8;
assign q[6519]= 16'h2da1;
assign q[6520]= 16'h2b59;
assign q[6521]= 16'h28fc;
assign q[6522]= 16'h2696;
assign q[6523]= 16'h2434;
assign q[6524]= 16'h21de;
assign q[6525]= 16'h1f9f;
assign q[6526]= 16'h1d7d;
assign q[6527]= 16'h1b81;
assign q[6528]= 16'h19ae;
assign q[6529]= 16'h180b;
assign q[6530]= 16'h169b;
assign q[6531]= 16'h1561;
assign q[6532]= 16'h145e;
assign q[6533]= 16'h1396;
assign q[6534]= 16'h1307;
assign q[6535]= 16'h12b4;
assign q[6536]= 16'h129c;
assign q[6537]= 16'h12be;
assign q[6538]= 16'h1319;
assign q[6539]= 16'h13ad;
assign q[6540]= 16'h1478;
assign q[6541]= 16'h1576;
assign q[6542]= 16'h16a7;
assign q[6543]= 16'h1806;
assign q[6544]= 16'h198f;
assign q[6545]= 16'h1b3f;
assign q[6546]= 16'h1d10;
assign q[6547]= 16'h1efc;
assign q[6548]= 16'h20fe;
assign q[6549]= 16'h230d;
assign q[6550]= 16'h2524;
assign q[6551]= 16'h2739;
assign q[6552]= 16'h2945;
assign q[6553]= 16'h2b3e;
assign q[6554]= 16'h2d1b;
assign q[6555]= 16'h2ed4;
assign q[6556]= 16'h305f;
assign q[6557]= 16'h31b4;
assign q[6558]= 16'h32c9;
assign q[6559]= 16'h3397;
assign q[6560]= 16'h3417;
assign q[6561]= 16'h3442;
assign q[6562]= 16'h3413;
assign q[6563]= 16'h3386;
assign q[6564]= 16'h3298;
assign q[6565]= 16'h3148;
assign q[6566]= 16'h2f96;
assign q[6567]= 16'h2d84;
assign q[6568]= 16'h2b17;
assign q[6569]= 16'h2853;
assign q[6570]= 16'h2540;
assign q[6571]= 16'h21e7;
assign q[6572]= 16'h1e52;
assign q[6573]= 16'h1a8e;
assign q[6574]= 16'h16a7;
assign q[6575]= 16'h12ac;
assign q[6576]= 16'heab;
assign q[6577]= 16'hab4;
assign q[6578]= 16'h6d6;
assign q[6579]= 16'h31f;
assign q[6580]= 16'hff9e;
assign q[6581]= 16'hfc5e;
assign q[6582]= 16'hf96a;
assign q[6583]= 16'hf6cd;
assign q[6584]= 16'hf48c;
assign q[6585]= 16'hf2ab;
assign q[6586]= 16'hf12e;
assign q[6587]= 16'hf011;
assign q[6588]= 16'hef51;
assign q[6589]= 16'heee8;
assign q[6590]= 16'heecb;
assign q[6591]= 16'heef0;
assign q[6592]= 16'hef48;
assign q[6593]= 16'hefc6;
assign q[6594]= 16'hf059;
assign q[6595]= 16'hf0f3;
assign q[6596]= 16'hf183;
assign q[6597]= 16'hf1fd;
assign q[6598]= 16'hf253;
assign q[6599]= 16'hf27c;
assign q[6600]= 16'hf271;
assign q[6601]= 16'hf22f;
assign q[6602]= 16'hf1b5;
assign q[6603]= 16'hf108;
assign q[6604]= 16'hf030;
assign q[6605]= 16'hef37;
assign q[6606]= 16'hee2e;
assign q[6607]= 16'hed24;
assign q[6608]= 16'hec2f;
assign q[6609]= 16'heb63;
assign q[6610]= 16'head6;
assign q[6611]= 16'hea9d;
assign q[6612]= 16'heacc;
assign q[6613]= 16'heb74;
assign q[6614]= 16'heca3;
assign q[6615]= 16'hee62;
assign q[6616]= 16'hf0b7;
assign q[6617]= 16'hf3a0;
assign q[6618]= 16'hf716;
assign q[6619]= 16'hfb0e;
assign q[6620]= 16'hff74;
assign q[6621]= 16'h430;
assign q[6622]= 16'h926;
assign q[6623]= 16'he35;
assign q[6624]= 16'h1339;
assign q[6625]= 16'h180d;
assign q[6626]= 16'h1c8b;
assign q[6627]= 16'h208e;
assign q[6628]= 16'h23f6;
assign q[6629]= 16'h26a3;
assign q[6630]= 16'h287e;
assign q[6631]= 16'h2974;
assign q[6632]= 16'h297b;
assign q[6633]= 16'h2890;
assign q[6634]= 16'h26ba;
assign q[6635]= 16'h2405;
assign q[6636]= 16'h208b;
assign q[6637]= 16'h1c68;
assign q[6638]= 16'h17c2;
assign q[6639]= 16'h12c4;
assign q[6640]= 16'hd9c;
assign q[6641]= 16'h87c;
assign q[6642]= 16'h393;
assign q[6643]= 16'hff14;
assign q[6644]= 16'hfb29;
assign q[6645]= 16'hf7fb;
assign q[6646]= 16'hf5a9;
assign q[6647]= 16'hf44e;
assign q[6648]= 16'hf3f8;
assign q[6649]= 16'hf4ac;
assign q[6650]= 16'hf667;
assign q[6651]= 16'hf917;
assign q[6652]= 16'hfca4;
assign q[6653]= 16'hea;
assign q[6654]= 16'h5c1;
assign q[6655]= 16'haf6;
assign q[6656]= 16'h1054;
assign q[6657]= 16'h15a4;
assign q[6658]= 16'h1aac;
assign q[6659]= 16'h1f36;
assign q[6660]= 16'h230f;
assign q[6661]= 16'h2609;
assign q[6662]= 16'h2801;
assign q[6663]= 16'h28da;
assign q[6664]= 16'h2882;
assign q[6665]= 16'h26f5;
assign q[6666]= 16'h2436;
assign q[6667]= 16'h2057;
assign q[6668]= 16'h1b75;
assign q[6669]= 16'h15b5;
assign q[6670]= 16'hf45;
assign q[6671]= 16'h85c;
assign q[6672]= 16'h134;
assign q[6673]= 16'hfa0b;
assign q[6674]= 16'hf31d;
assign q[6675]= 16'heca8;
assign q[6676]= 16'he6e2;
assign q[6677]= 16'he200;
assign q[6678]= 16'hde2a;
assign q[6679]= 16'hdb82;
assign q[6680]= 16'hda1e;
assign q[6681]= 16'hda09;
assign q[6682]= 16'hdb42;
assign q[6683]= 16'hddbe;
assign q[6684]= 16'he165;
assign q[6685]= 16'he616;
assign q[6686]= 16'heba7;
assign q[6687]= 16'hf1e8;
assign q[6688]= 16'hf8a2;
assign q[6689]= 16'hff9d;
assign q[6690]= 16'h69d;
assign q[6691]= 16'hd6a;
assign q[6692]= 16'h13ce;
assign q[6693]= 16'h1997;
assign q[6694]= 16'h1e99;
assign q[6695]= 16'h22b3;
assign q[6696]= 16'h25c9;
assign q[6697]= 16'h27ca;
assign q[6698]= 16'h28b0;
assign q[6699]= 16'h287d;
assign q[6700]= 16'h273e;
assign q[6701]= 16'h2507;
assign q[6702]= 16'h21f3;
assign q[6703]= 16'h1e25;
assign q[6704]= 16'h19c5;
assign q[6705]= 16'h14fb;
assign q[6706]= 16'hff5;
assign q[6707]= 16'hadd;
assign q[6708]= 16'h5de;
assign q[6709]= 16'h11f;
assign q[6710]= 16'hfcc4;
assign q[6711]= 16'hf8e9;
assign q[6712]= 16'hf5a9;
assign q[6713]= 16'hf314;
assign q[6714]= 16'hf136;
assign q[6715]= 16'hf015;
assign q[6716]= 16'hefaf;
assign q[6717]= 16'heffe;
assign q[6718]= 16'hf0f4;
assign q[6719]= 16'hf283;
assign q[6720]= 16'hf495;
assign q[6721]= 16'hf715;
assign q[6722]= 16'hf9eb;
assign q[6723]= 16'hfcfe;
assign q[6724]= 16'h35;
assign q[6725]= 16'h379;
assign q[6726]= 16'h6b4;
assign q[6727]= 16'h9d2;
assign q[6728]= 16'hcc0;
assign q[6729]= 16'hf6f;
assign q[6730]= 16'h11d3;
assign q[6731]= 16'h13e2;
assign q[6732]= 16'h1595;
assign q[6733]= 16'h16e6;
assign q[6734]= 16'h17d5;
assign q[6735]= 16'h1860;
assign q[6736]= 16'h1888;
assign q[6737]= 16'h1851;
assign q[6738]= 16'h17bd;
assign q[6739]= 16'h16d3;
assign q[6740]= 16'h1599;
assign q[6741]= 16'h1415;
assign q[6742]= 16'h124e;
assign q[6743]= 16'h104d;
assign q[6744]= 16'he1c;
assign q[6745]= 16'hbc2;
assign q[6746]= 16'h94c;
assign q[6747]= 16'h6c3;
assign q[6748]= 16'h433;
assign q[6749]= 16'h1a9;
assign q[6750]= 16'hff31;
assign q[6751]= 16'hfcd7;
assign q[6752]= 16'hfaa7;
assign q[6753]= 16'hf8ae;
assign q[6754]= 16'hf6f8;
assign q[6755]= 16'hf58f;
assign q[6756]= 16'hf47c;
assign q[6757]= 16'hf3c6;
assign q[6758]= 16'hf372;
assign q[6759]= 16'hf383;
assign q[6760]= 16'hf3f9;
assign q[6761]= 16'hf4d0;
assign q[6762]= 16'hf602;
assign q[6763]= 16'hf786;
assign q[6764]= 16'hf950;
assign q[6765]= 16'hfb52;
assign q[6766]= 16'hfd7a;
assign q[6767]= 16'hffb5;
assign q[6768]= 16'h1ef;
assign q[6769]= 16'h416;
assign q[6770]= 16'h612;
assign q[6771]= 16'h7d1;
assign q[6772]= 16'h93f;
assign q[6773]= 16'ha4b;
assign q[6774]= 16'hae8;
assign q[6775]= 16'hb0a;
assign q[6776]= 16'haa8;
assign q[6777]= 16'h9c0;
assign q[6778]= 16'h851;
assign q[6779]= 16'h65f;
assign q[6780]= 16'h3f0;
assign q[6781]= 16'h110;
assign q[6782]= 16'hfdcf;
assign q[6783]= 16'hfa3b;
assign q[6784]= 16'hf669;
assign q[6785]= 16'hf26e;
assign q[6786]= 16'hee5f;
assign q[6787]= 16'hea54;
assign q[6788]= 16'he662;
assign q[6789]= 16'he29f;
assign q[6790]= 16'hdf1f;
assign q[6791]= 16'hdbf4;
assign q[6792]= 16'hd92e;
assign q[6793]= 16'hd6db;
assign q[6794]= 16'hd507;
assign q[6795]= 16'hd3b8;
assign q[6796]= 16'hd2f6;
assign q[6797]= 16'hd2c2;
assign q[6798]= 16'hd31d;
assign q[6799]= 16'hd406;
assign q[6800]= 16'hd577;
assign q[6801]= 16'hd76c;
assign q[6802]= 16'hd9db;
assign q[6803]= 16'hdcbe;
assign q[6804]= 16'he008;
assign q[6805]= 16'he3af;
assign q[6806]= 16'he7a7;
assign q[6807]= 16'hebe3;
assign q[6808]= 16'hf056;
assign q[6809]= 16'hf4f3;
assign q[6810]= 16'hf9ab;
assign q[6811]= 16'hfe70;
assign q[6812]= 16'h333;
assign q[6813]= 16'h7e6;
assign q[6814]= 16'hc79;
assign q[6815]= 16'h10df;
assign q[6816]= 16'h1508;
assign q[6817]= 16'h18e7;
assign q[6818]= 16'h1c6e;
assign q[6819]= 16'h1f92;
assign q[6820]= 16'h2248;
assign q[6821]= 16'h2486;
assign q[6822]= 16'h2647;
assign q[6823]= 16'h2786;
assign q[6824]= 16'h2841;
assign q[6825]= 16'h2879;
assign q[6826]= 16'h2832;
assign q[6827]= 16'h2775;
assign q[6828]= 16'h264a;
assign q[6829]= 16'h24c0;
assign q[6830]= 16'h22e6;
assign q[6831]= 16'h20ce;
assign q[6832]= 16'h1e8c;
assign q[6833]= 16'h1c33;
assign q[6834]= 16'h19da;
assign q[6835]= 16'h1795;
assign q[6836]= 16'h1576;
assign q[6837]= 16'h1390;
assign q[6838]= 16'h11f0;
assign q[6839]= 16'h10a3;
assign q[6840]= 16'hfb0;
assign q[6841]= 16'hf19;
assign q[6842]= 16'hedf;
assign q[6843]= 16'hefa;
assign q[6844]= 16'hf61;
assign q[6845]= 16'h1005;
assign q[6846]= 16'h10d3;
assign q[6847]= 16'h11b7;
assign q[6848]= 16'h1298;
assign q[6849]= 16'h135e;
assign q[6850]= 16'h13ef;
assign q[6851]= 16'h1433;
assign q[6852]= 16'h1415;
assign q[6853]= 16'h1380;
assign q[6854]= 16'h1266;
assign q[6855]= 16'h10bb;
assign q[6856]= 16'he7b;
assign q[6857]= 16'hba7;
assign q[6858]= 16'h845;
assign q[6859]= 16'h464;
assign q[6860]= 16'h17;
assign q[6861]= 16'hfb77;
assign q[6862]= 16'hf6a1;
assign q[6863]= 16'hf1b7;
assign q[6864]= 16'hecdd;
assign q[6865]= 16'he83a;
assign q[6866]= 16'he3f3;
assign q[6867]= 16'he02e;
assign q[6868]= 16'hdd0d;
assign q[6869]= 16'hdaad;
assign q[6870]= 16'hd928;
assign q[6871]= 16'hd891;
assign q[6872]= 16'hd8f5;
assign q[6873]= 16'hda57;
assign q[6874]= 16'hdcb4;
assign q[6875]= 16'he002;
assign q[6876]= 16'he42d;
assign q[6877]= 16'he91b;
assign q[6878]= 16'heeac;
assign q[6879]= 16'hf4bb;
assign q[6880]= 16'hfb1d;
assign q[6881]= 16'h1a6;
assign q[6882]= 16'h82a;
assign q[6883]= 16'he7a;
assign q[6884]= 16'h146a;
assign q[6885]= 16'h19d3;
assign q[6886]= 16'h1e8f;
assign q[6887]= 16'h2280;
assign q[6888]= 16'h258d;
assign q[6889]= 16'h27a5;
assign q[6890]= 16'h28bf;
assign q[6891]= 16'h28d7;
assign q[6892]= 16'h27f4;
assign q[6893]= 16'h2621;
assign q[6894]= 16'h2371;
assign q[6895]= 16'h1ffc;
assign q[6896]= 16'h1bdf;
assign q[6897]= 16'h173a;
assign q[6898]= 16'h1230;
assign q[6899]= 16'hce4;
assign q[6900]= 16'h779;
assign q[6901]= 16'h210;
assign q[6902]= 16'hfcc8;
assign q[6903]= 16'hf7bc;
assign q[6904]= 16'hf302;
assign q[6905]= 16'heeac;
assign q[6906]= 16'heac8;
assign q[6907]= 16'he75c;
assign q[6908]= 16'he46b;
assign q[6909]= 16'he1f1;
assign q[6910]= 16'hdfe8;
assign q[6911]= 16'hde44;
assign q[6912]= 16'hdcf7;
assign q[6913]= 16'hdbf2;
assign q[6914]= 16'hdb23;
assign q[6915]= 16'hda79;
assign q[6916]= 16'hd9e4;
assign q[6917]= 16'hd954;
assign q[6918]= 16'hd8bc;
assign q[6919]= 16'hd812;
assign q[6920]= 16'hd750;
assign q[6921]= 16'hd672;
assign q[6922]= 16'hd57a;
assign q[6923]= 16'hd46b;
assign q[6924]= 16'hd34c;
assign q[6925]= 16'hd229;
assign q[6926]= 16'hd10e;
assign q[6927]= 16'hd009;
assign q[6928]= 16'hcf2b;
assign q[6929]= 16'hce84;
assign q[6930]= 16'hce23;
assign q[6931]= 16'hce16;
assign q[6932]= 16'hce6a;
assign q[6933]= 16'hcf2a;
assign q[6934]= 16'hd05c;
assign q[6935]= 16'hd204;
assign q[6936]= 16'hd422;
assign q[6937]= 16'hd6b2;
assign q[6938]= 16'hd9ad;
assign q[6939]= 16'hdd08;
assign q[6940]= 16'he0b5;
assign q[6941]= 16'he4a3;
assign q[6942]= 16'he8bf;
assign q[6943]= 16'hecf5;
assign q[6944]= 16'hf12e;
assign q[6945]= 16'hf556;
assign q[6946]= 16'hf957;
assign q[6947]= 16'hfd1d;
assign q[6948]= 16'h93;
assign q[6949]= 16'h3ac;
assign q[6950]= 16'h659;
assign q[6951]= 16'h88f;
assign q[6952]= 16'ha46;
assign q[6953]= 16'hb7b;
assign q[6954]= 16'hc2b;
assign q[6955]= 16'hc5a;
assign q[6956]= 16'hc0c;
assign q[6957]= 16'hb49;
assign q[6958]= 16'ha1b;
assign q[6959]= 16'h88f;
assign q[6960]= 16'h6b3;
assign q[6961]= 16'h494;
assign q[6962]= 16'h243;
assign q[6963]= 16'hffcf;
assign q[6964]= 16'hfd47;
assign q[6965]= 16'hfaba;
assign q[6966]= 16'hf835;
assign q[6967]= 16'hf5c6;
assign q[6968]= 16'hf379;
assign q[6969]= 16'hf158;
assign q[6970]= 16'hef6b;
assign q[6971]= 16'hedba;
assign q[6972]= 16'hec4c;
assign q[6973]= 16'heb26;
assign q[6974]= 16'hea4b;
assign q[6975]= 16'he9be;
assign q[6976]= 16'he982;
assign q[6977]= 16'he998;
assign q[6978]= 16'hea00;
assign q[6979]= 16'heaba;
assign q[6980]= 16'hebc5;
assign q[6981]= 16'hed21;
assign q[6982]= 16'heecc;
assign q[6983]= 16'hf0c4;
assign q[6984]= 16'hf304;
assign q[6985]= 16'hf58b;
assign q[6986]= 16'hf853;
assign q[6987]= 16'hfb57;
assign q[6988]= 16'hfe91;
assign q[6989]= 16'h1f9;
assign q[6990]= 16'h589;
assign q[6991]= 16'h936;
assign q[6992]= 16'hcf7;
assign q[6993]= 16'h10c2;
assign q[6994]= 16'h148b;
assign q[6995]= 16'h1847;
assign q[6996]= 16'h1beb;
assign q[6997]= 16'h1f6a;
assign q[6998]= 16'h22bb;
assign q[6999]= 16'h25d2;
assign q[7000]= 16'h28a6;
assign q[7001]= 16'h2b2e;
assign q[7002]= 16'h2d64;
assign q[7003]= 16'h2f43;
assign q[7004]= 16'h30c5;
assign q[7005]= 16'h31ea;
assign q[7006]= 16'h32b1;
assign q[7007]= 16'h331b;
assign q[7008]= 16'h332b;
assign q[7009]= 16'h32e4;
assign q[7010]= 16'h324d;
assign q[7011]= 16'h316a;
assign q[7012]= 16'h3043;
assign q[7013]= 16'h2edd;
assign q[7014]= 16'h2d40;
assign q[7015]= 16'h2b71;
assign q[7016]= 16'h2975;
assign q[7017]= 16'h2751;
assign q[7018]= 16'h2508;
assign q[7019]= 16'h229c;
assign q[7020]= 16'h200f;
assign q[7021]= 16'h1d5f;
assign q[7022]= 16'h1a8d;
assign q[7023]= 16'h1796;
assign q[7024]= 16'h1478;
assign q[7025]= 16'h1133;
assign q[7026]= 16'hdc3;
assign q[7027]= 16'ha28;
assign q[7028]= 16'h663;
assign q[7029]= 16'h276;
assign q[7030]= 16'hfe64;
assign q[7031]= 16'hfa32;
assign q[7032]= 16'hf5ea;
assign q[7033]= 16'hf195;
assign q[7034]= 16'hed42;
assign q[7035]= 16'he8fd;
assign q[7036]= 16'he4da;
assign q[7037]= 16'he0ea;
assign q[7038]= 16'hdd42;
assign q[7039]= 16'hd9f5;
assign q[7040]= 16'hd718;
assign q[7041]= 16'hd4be;
assign q[7042]= 16'hd2f9;
assign q[7043]= 16'hd1d9;
assign q[7044]= 16'hd16b;
assign q[7045]= 16'hd1b9;
assign q[7046]= 16'hd2c8;
assign q[7047]= 16'hd49b;
assign q[7048]= 16'hd72d;
assign q[7049]= 16'hda76;
assign q[7050]= 16'hde6b;
assign q[7051]= 16'he2fb;
assign q[7052]= 16'he810;
assign q[7053]= 16'hed91;
assign q[7054]= 16'hf364;
assign q[7055]= 16'hf96a;
assign q[7056]= 16'hff84;
assign q[7057]= 16'h592;
assign q[7058]= 16'hb75;
assign q[7059]= 16'h1110;
assign q[7060]= 16'h1646;
assign q[7061]= 16'h1aff;
assign q[7062]= 16'h1f25;
assign q[7063]= 16'h22a8;
assign q[7064]= 16'h257b;
assign q[7065]= 16'h2799;
assign q[7066]= 16'h28ff;
assign q[7067]= 16'h29b0;
assign q[7068]= 16'h29b6;
assign q[7069]= 16'h291d;
assign q[7070]= 16'h27f5;
assign q[7071]= 16'h2654;
assign q[7072]= 16'h2451;
assign q[7073]= 16'h2204;
assign q[7074]= 16'h1f88;
assign q[7075]= 16'h1cf7;
assign q[7076]= 16'h1a6b;
assign q[7077]= 16'h17fd;
assign q[7078]= 16'h15c2;
assign q[7079]= 16'h13d0;
assign q[7080]= 16'h1237;
assign q[7081]= 16'h1104;
assign q[7082]= 16'h1041;
assign q[7083]= 16'hff3;
assign q[7084]= 16'h101d;
assign q[7085]= 16'h10be;
assign q[7086]= 16'h11cf;
assign q[7087]= 16'h1349;
assign q[7088]= 16'h1521;
assign q[7089]= 16'h174a;
assign q[7090]= 16'h19b6;
assign q[7091]= 16'h1c55;
assign q[7092]= 16'h1f15;
assign q[7093]= 16'h21e7;
assign q[7094]= 16'h24ba;
assign q[7095]= 16'h277e;
assign q[7096]= 16'h2a24;
assign q[7097]= 16'h2c9d;
assign q[7098]= 16'h2ede;
assign q[7099]= 16'h30dc;
assign q[7100]= 16'h328e;
assign q[7101]= 16'h33eb;
assign q[7102]= 16'h34ee;
assign q[7103]= 16'h3592;
assign q[7104]= 16'h35d4;
assign q[7105]= 16'h35b3;
assign q[7106]= 16'h352e;
assign q[7107]= 16'h3446;
assign q[7108]= 16'h32fd;
assign q[7109]= 16'h3157;
assign q[7110]= 16'h2f57;
assign q[7111]= 16'h2d03;
assign q[7112]= 16'h2a61;
assign q[7113]= 16'h2778;
assign q[7114]= 16'h2450;
assign q[7115]= 16'h20f2;
assign q[7116]= 16'h1d67;
assign q[7117]= 16'h19ba;
assign q[7118]= 16'h15f5;
assign q[7119]= 16'h1226;
assign q[7120]= 16'he56;
assign q[7121]= 16'ha93;
assign q[7122]= 16'h6e9;
assign q[7123]= 16'h362;
assign q[7124]= 16'hb;
assign q[7125]= 16'hfcee;
assign q[7126]= 16'hfa12;
assign q[7127]= 16'hf780;
assign q[7128]= 16'hf53e;
assign q[7129]= 16'hf34f;
assign q[7130]= 16'hf1b5;
assign q[7131]= 16'hf071;
assign q[7132]= 16'hef7f;
assign q[7133]= 16'heedb;
assign q[7134]= 16'hee7e;
assign q[7135]= 16'hee60;
assign q[7136]= 16'hee78;
assign q[7137]= 16'heeba;
assign q[7138]= 16'hef1a;
assign q[7139]= 16'hef8d;
assign q[7140]= 16'hf006;
assign q[7141]= 16'hf07b;
assign q[7142]= 16'hf0e1;
assign q[7143]= 16'hf130;
assign q[7144]= 16'hf162;
assign q[7145]= 16'hf172;
assign q[7146]= 16'hf15f;
assign q[7147]= 16'hf129;
assign q[7148]= 16'hf0d4;
assign q[7149]= 16'hf067;
assign q[7150]= 16'hefea;
assign q[7151]= 16'hef67;
assign q[7152]= 16'heeea;
assign q[7153]= 16'hee83;
assign q[7154]= 16'hee3d;
assign q[7155]= 16'hee29;
assign q[7156]= 16'hee53;
assign q[7157]= 16'heec8;
assign q[7158]= 16'hef93;
assign q[7159]= 16'hf0be;
assign q[7160]= 16'hf24e;
assign q[7161]= 16'hf446;
assign q[7162]= 16'hf6a7;
assign q[7163]= 16'hf96d;
assign q[7164]= 16'hfc91;
assign q[7165]= 16'h9;
assign q[7166]= 16'h3c9;
assign q[7167]= 16'h7c2;
assign q[7168]= 16'hbe2;
assign q[7169]= 16'h1015;
assign q[7170]= 16'h1449;
assign q[7171]= 16'h1868;
assign q[7172]= 16'h1c61;
assign q[7173]= 16'h2020;
assign q[7174]= 16'h2395;
assign q[7175]= 16'h26b2;
assign q[7176]= 16'h296c;
assign q[7177]= 16'h2bbb;
assign q[7178]= 16'h2d9b;
assign q[7179]= 16'h2f0a;
assign q[7180]= 16'h300b;
assign q[7181]= 16'h30a4;
assign q[7182]= 16'h30df;
assign q[7183]= 16'h30c6;
assign q[7184]= 16'h3069;
assign q[7185]= 16'h2fd6;
assign q[7186]= 16'h2f1d;
assign q[7187]= 16'h2e50;
assign q[7188]= 16'h2d7e;
assign q[7189]= 16'h2cb6;
assign q[7190]= 16'h2c06;
assign q[7191]= 16'h2b79;
assign q[7192]= 16'h2b15;
assign q[7193]= 16'h2ae2;
assign q[7194]= 16'h2ae0;
assign q[7195]= 16'h2b0f;
assign q[7196]= 16'h2b69;
assign q[7197]= 16'h2be8;
assign q[7198]= 16'h2c82;
assign q[7199]= 16'h2d2a;
assign q[7200]= 16'h2dd3;
assign q[7201]= 16'h2e6e;
assign q[7202]= 16'h2eee;
assign q[7203]= 16'h2f43;
assign q[7204]= 16'h2f61;
assign q[7205]= 16'h2f3c;
assign q[7206]= 16'h2ecc;
assign q[7207]= 16'h2e0b;
assign q[7208]= 16'h2cf5;
assign q[7209]= 16'h2b8d;
assign q[7210]= 16'h29d4;
assign q[7211]= 16'h27d4;
assign q[7212]= 16'h2598;
assign q[7213]= 16'h232c;
assign q[7214]= 16'h20a1;
assign q[7215]= 16'h1e0a;
assign q[7216]= 16'h1b79;
assign q[7217]= 16'h1903;
assign q[7218]= 16'h16bb;
assign q[7219]= 16'h14b3;
assign q[7220]= 16'h12fd;
assign q[7221]= 16'h11a7;
assign q[7222]= 16'h10bb;
assign q[7223]= 16'h1043;
assign q[7224]= 16'h1042;
assign q[7225]= 16'h10b8;
assign q[7226]= 16'h11a0;
assign q[7227]= 16'h12f3;
assign q[7228]= 16'h14a5;
assign q[7229]= 16'h16a5;
assign q[7230]= 16'h18e3;
assign q[7231]= 16'h1b49;
assign q[7232]= 16'h1dc1;
assign q[7233]= 16'h2035;
assign q[7234]= 16'h228e;
assign q[7235]= 16'h24b7;
assign q[7236]= 16'h269c;
assign q[7237]= 16'h282b;
assign q[7238]= 16'h2956;
assign q[7239]= 16'h2a12;
assign q[7240]= 16'h2a59;
assign q[7241]= 16'h2a28;
assign q[7242]= 16'h2981;
assign q[7243]= 16'h286b;
assign q[7244]= 16'h26ef;
assign q[7245]= 16'h251d;
assign q[7246]= 16'h2304;
assign q[7247]= 16'h20b8;
assign q[7248]= 16'h1e50;
assign q[7249]= 16'h1be1;
assign q[7250]= 16'h1983;
assign q[7251]= 16'h174a;
assign q[7252]= 16'h154d;
assign q[7253]= 16'h139e;
assign q[7254]= 16'h124b;
assign q[7255]= 16'h1161;
assign q[7256]= 16'h10e9;
assign q[7257]= 16'h10e7;
assign q[7258]= 16'h115a;
assign q[7259]= 16'h123e;
assign q[7260]= 16'h138b;
assign q[7261]= 16'h1534;
assign q[7262]= 16'h172a;
assign q[7263]= 16'h195b;
assign q[7264]= 16'h1bb2;
assign q[7265]= 16'h1e1a;
assign q[7266]= 16'h207d;
assign q[7267]= 16'h22c5;
assign q[7268]= 16'h24dd;
assign q[7269]= 16'h26b3;
assign q[7270]= 16'h2835;
assign q[7271]= 16'h2957;
assign q[7272]= 16'h2a0e;
assign q[7273]= 16'h2a54;
assign q[7274]= 16'h2a27;
assign q[7275]= 16'h2989;
assign q[7276]= 16'h287f;
assign q[7277]= 16'h2712;
assign q[7278]= 16'h254f;
assign q[7279]= 16'h2345;
assign q[7280]= 16'h2106;
assign q[7281]= 16'h1ea2;
assign q[7282]= 16'h1c2f;
assign q[7283]= 16'h19c0;
assign q[7284]= 16'h1766;
assign q[7285]= 16'h1532;
assign q[7286]= 16'h1335;
assign q[7287]= 16'h117a;
assign q[7288]= 16'h1009;
assign q[7289]= 16'hee9;
assign q[7290]= 16'he1c;
assign q[7291]= 16'hda0;
assign q[7292]= 16'hd6e;
assign q[7293]= 16'hd7f;
assign q[7294]= 16'hdc7;
assign q[7295]= 16'he36;
assign q[7296]= 16'hebc;
assign q[7297]= 16'hf47;
assign q[7298]= 16'hfc4;
assign q[7299]= 16'h1020;
assign q[7300]= 16'h1048;
assign q[7301]= 16'h102c;
assign q[7302]= 16'hfbc;
assign q[7303]= 16'heed;
assign q[7304]= 16'hdb5;
assign q[7305]= 16'hc0d;
assign q[7306]= 16'h9f5;
assign q[7307]= 16'h76c;
assign q[7308]= 16'h47a;
assign q[7309]= 16'h126;
assign q[7310]= 16'hfd7f;
assign q[7311]= 16'hf990;
assign q[7312]= 16'hf56d;
assign q[7313]= 16'hf12a;
assign q[7314]= 16'hecda;
assign q[7315]= 16'he893;
assign q[7316]= 16'he469;
assign q[7317]= 16'he070;
assign q[7318]= 16'hdcba;
assign q[7319]= 16'hd958;
assign q[7320]= 16'hd656;
assign q[7321]= 16'hd3bf;
assign q[7322]= 16'hd199;
assign q[7323]= 16'hcfe9;
assign q[7324]= 16'hcead;
assign q[7325]= 16'hcde3;
assign q[7326]= 16'hcd84;
assign q[7327]= 16'hcd87;
assign q[7328]= 16'hcde0;
assign q[7329]= 16'hce82;
assign q[7330]= 16'hcf5f;
assign q[7331]= 16'hd069;
assign q[7332]= 16'hd191;
assign q[7333]= 16'hd2c9;
assign q[7334]= 16'hd406;
assign q[7335]= 16'hd53e;
assign q[7336]= 16'hd66a;
assign q[7337]= 16'hd784;
assign q[7338]= 16'hd88c;
assign q[7339]= 16'hd981;
assign q[7340]= 16'hda68;
assign q[7341]= 16'hdb47;
assign q[7342]= 16'hdc27;
assign q[7343]= 16'hdd12;
assign q[7344]= 16'hde13;
assign q[7345]= 16'hdf37;
assign q[7346]= 16'he088;
assign q[7347]= 16'he211;
assign q[7348]= 16'he3db;
assign q[7349]= 16'he5eb;
assign q[7350]= 16'he847;
assign q[7351]= 16'heaed;
assign q[7352]= 16'hedda;
assign q[7353]= 16'hf106;
assign q[7354]= 16'hf466;
assign q[7355]= 16'hf7ec;
assign q[7356]= 16'hfb85;
assign q[7357]= 16'hff1b;
assign q[7358]= 16'h297;
assign q[7359]= 16'h5e2;
assign q[7360]= 16'h8e2;
assign q[7361]= 16'hb7e;
assign q[7362]= 16'hd9f;
assign q[7363]= 16'hf30;
assign q[7364]= 16'h101f;
assign q[7365]= 16'h1060;
assign q[7366]= 16'hfea;
assign q[7367]= 16'heba;
assign q[7368]= 16'hcd2;
assign q[7369]= 16'ha3c;
assign q[7370]= 16'h705;
assign q[7371]= 16'h342;
assign q[7372]= 16'hff0e;
assign q[7373]= 16'hfa84;
assign q[7374]= 16'hf5c7;
assign q[7375]= 16'hf0fb;
assign q[7376]= 16'hec47;
assign q[7377]= 16'he7cf;
assign q[7378]= 16'he3ba;
assign q[7379]= 16'he02b;
assign q[7380]= 16'hdd41;
assign q[7381]= 16'hdb18;
assign q[7382]= 16'hd9c6;
assign q[7383]= 16'hd95a;
assign q[7384]= 16'hd9de;
assign q[7385]= 16'hdb54;
assign q[7386]= 16'hddb7;
assign q[7387]= 16'he0fa;
assign q[7388]= 16'he50b;
assign q[7389]= 16'he9d1;
assign q[7390]= 16'hef2e;
assign q[7391]= 16'hf4fe;
assign q[7392]= 16'hfb1b;
assign q[7393]= 16'h15c;
assign q[7394]= 16'h799;
assign q[7395]= 16'hda9;
assign q[7396]= 16'h1363;
assign q[7397]= 16'h18a4;
assign q[7398]= 16'h1d4b;
assign q[7399]= 16'h213a;
assign q[7400]= 16'h245b;
assign q[7401]= 16'h269c;
assign q[7402]= 16'h27f4;
assign q[7403]= 16'h285d;
assign q[7404]= 16'h27d9;
assign q[7405]= 16'h266f;
assign q[7406]= 16'h242e;
assign q[7407]= 16'h2128;
assign q[7408]= 16'h1d72;
assign q[7409]= 16'h1927;
assign q[7410]= 16'h1462;
assign q[7411]= 16'hf42;
assign q[7412]= 16'h9e4;
assign q[7413]= 16'h467;
assign q[7414]= 16'hfee8;
assign q[7415]= 16'hf980;
assign q[7416]= 16'hf448;
assign q[7417]= 16'hef56;
assign q[7418]= 16'heabb;
assign q[7419]= 16'he687;
assign q[7420]= 16'he2c3;
assign q[7421]= 16'hdf77;
assign q[7422]= 16'hdca6;
assign q[7423]= 16'hda52;
assign q[7424]= 16'hd877;
assign q[7425]= 16'hd711;
assign q[7426]= 16'hd619;
assign q[7427]= 16'hd588;
assign q[7428]= 16'hd553;
assign q[7429]= 16'hd571;
assign q[7430]= 16'hd5d7;
assign q[7431]= 16'hd67c;
assign q[7432]= 16'hd756;
assign q[7433]= 16'hd85b;
assign q[7434]= 16'hd985;
assign q[7435]= 16'hdacc;
assign q[7436]= 16'hdc29;
assign q[7437]= 16'hdd98;
assign q[7438]= 16'hdf13;
assign q[7439]= 16'he097;
assign q[7440]= 16'he221;
assign q[7441]= 16'he3ad;
assign q[7442]= 16'he53a;
assign q[7443]= 16'he6c5;
assign q[7444]= 16'he84b;
assign q[7445]= 16'he9ca;
assign q[7446]= 16'heb3f;
assign q[7447]= 16'heca8;
assign q[7448]= 16'hee00;
assign q[7449]= 16'hef45;
assign q[7450]= 16'hf073;
assign q[7451]= 16'hf186;
assign q[7452]= 16'hf27b;
assign q[7453]= 16'hf34e;
assign q[7454]= 16'hf3fc;
assign q[7455]= 16'hf483;
assign q[7456]= 16'hf4df;
assign q[7457]= 16'hf511;
assign q[7458]= 16'hf518;
assign q[7459]= 16'hf4f3;
assign q[7460]= 16'hf4a5;
assign q[7461]= 16'hf431;
assign q[7462]= 16'hf39a;
assign q[7463]= 16'hf2e5;
assign q[7464]= 16'hf218;
assign q[7465]= 16'hf139;
assign q[7466]= 16'hf052;
assign q[7467]= 16'hef69;
assign q[7468]= 16'hee88;
assign q[7469]= 16'hedb8;
assign q[7470]= 16'hed03;
assign q[7471]= 16'hec73;
assign q[7472]= 16'hec11;
assign q[7473]= 16'hebe5;
assign q[7474]= 16'hebf8;
assign q[7475]= 16'hec51;
assign q[7476]= 16'hecf6;
assign q[7477]= 16'hedec;
assign q[7478]= 16'hef37;
assign q[7479]= 16'hf0d7;
assign q[7480]= 16'hf2ce;
assign q[7481]= 16'hf51a;
assign q[7482]= 16'hf7b6;
assign q[7483]= 16'hfa9f;
assign q[7484]= 16'hfdcc;
assign q[7485]= 16'h135;
assign q[7486]= 16'h4d1;
assign q[7487]= 16'h893;
assign q[7488]= 16'hc71;
assign q[7489]= 16'h105b;
assign q[7490]= 16'h1445;
assign q[7491]= 16'h1822;
assign q[7492]= 16'h1be2;
assign q[7493]= 16'h1f7a;
assign q[7494]= 16'h22de;
assign q[7495]= 16'h2601;
assign q[7496]= 16'h28da;
assign q[7497]= 16'h2b61;
assign q[7498]= 16'h2d90;
assign q[7499]= 16'h2f62;
assign q[7500]= 16'h30d5;
assign q[7501]= 16'h31e7;
assign q[7502]= 16'h329a;
assign q[7503]= 16'h32f1;
assign q[7504]= 16'h32ef;
assign q[7505]= 16'h329b;
assign q[7506]= 16'h31fa;
assign q[7507]= 16'h3112;
assign q[7508]= 16'h2fec;
assign q[7509]= 16'h2e8d;
assign q[7510]= 16'h2cfd;
assign q[7511]= 16'h2b3f;
assign q[7512]= 16'h295a;
assign q[7513]= 16'h274f;
assign q[7514]= 16'h2522;
assign q[7515]= 16'h22d3;
assign q[7516]= 16'h2062;
assign q[7517]= 16'h1dcc;
assign q[7518]= 16'h1b11;
assign q[7519]= 16'h182b;
assign q[7520]= 16'h151a;
assign q[7521]= 16'h11d9;
assign q[7522]= 16'he67;
assign q[7523]= 16'hac1;
assign q[7524]= 16'h6ea;
assign q[7525]= 16'h2e2;
assign q[7526]= 16'hfeb0;
assign q[7527]= 16'hfa58;
assign q[7528]= 16'hf5e5;
assign q[7529]= 16'hf162;
assign q[7530]= 16'hece0;
assign q[7531]= 16'he86e;
assign q[7532]= 16'he421;
assign q[7533]= 16'he00c;
assign q[7534]= 16'hdc45;
assign q[7535]= 16'hd8e3;
assign q[7536]= 16'hd5fb;
assign q[7537]= 16'hd3a3;
assign q[7538]= 16'hd1ec;
assign q[7539]= 16'hd0e8;
assign q[7540]= 16'hd0a3;
assign q[7541]= 16'hd127;
assign q[7542]= 16'hd279;
assign q[7543]= 16'hd498;
assign q[7544]= 16'hd77f;
assign q[7545]= 16'hdb24;
assign q[7546]= 16'hdf78;
assign q[7547]= 16'he465;
assign q[7548]= 16'he9d3;
assign q[7549]= 16'hefa5;
assign q[7550]= 16'hf5ba;
assign q[7551]= 16'hfbef;
assign q[7552]= 16'h220;
assign q[7553]= 16'h828;
assign q[7554]= 16'hde3;
assign q[7555]= 16'h132e;
assign q[7556]= 16'h17e6;
assign q[7557]= 16'h1bee;
assign q[7558]= 16'h1f2e;
assign q[7559]= 16'h218f;
assign q[7560]= 16'h2302;
assign q[7561]= 16'h237e;
assign q[7562]= 16'h22ff;
assign q[7563]= 16'h2186;
assign q[7564]= 16'h1f1c;
assign q[7565]= 16'h1bce;
assign q[7566]= 16'h17af;
assign q[7567]= 16'h12d6;
assign q[7568]= 16'hd5e;
assign q[7569]= 16'h765;
assign q[7570]= 16'h10d;
assign q[7571]= 16'hfa78;
assign q[7572]= 16'hf3c7;
assign q[7573]= 16'hed1d;
assign q[7574]= 16'he69b;
assign q[7575]= 16'he060;
assign q[7576]= 16'hda89;
assign q[7577]= 16'hd52f;
assign q[7578]= 16'hd06a;
assign q[7579]= 16'hcc4a;
assign q[7580]= 16'hc8de;
assign q[7581]= 16'hc62f;
assign q[7582]= 16'hc443;
assign q[7583]= 16'hc31c;
assign q[7584]= 16'hc2b8;
assign q[7585]= 16'hc30f;
assign q[7586]= 16'hc419;
assign q[7587]= 16'hc5ca;
assign q[7588]= 16'hc814;
assign q[7589]= 16'hcae5;
assign q[7590]= 16'hce2b;
assign q[7591]= 16'hd1d4;
assign q[7592]= 16'hd5cb;
assign q[7593]= 16'hd9fd;
assign q[7594]= 16'hde54;
assign q[7595]= 16'he2be;
assign q[7596]= 16'he728;
assign q[7597]= 16'heb7e;
assign q[7598]= 16'hefb1;
assign q[7599]= 16'hf3b0;
assign q[7600]= 16'hf76d;
assign q[7601]= 16'hfada;
assign q[7602]= 16'hfded;
assign q[7603]= 16'h9a;
assign q[7604]= 16'h2dc;
assign q[7605]= 16'h4a9;
assign q[7606]= 16'h5fe;
assign q[7607]= 16'h6d6;
assign q[7608]= 16'h730;
assign q[7609]= 16'h70b;
assign q[7610]= 16'h669;
assign q[7611]= 16'h54b;
assign q[7612]= 16'h3b6;
assign q[7613]= 16'h1b0;
assign q[7614]= 16'hff41;
assign q[7615]= 16'hfc70;
assign q[7616]= 16'hf946;
assign q[7617]= 16'hf5d1;
assign q[7618]= 16'hf21c;
assign q[7619]= 16'hee34;
assign q[7620]= 16'hea2a;
assign q[7621]= 16'he60b;
assign q[7622]= 16'he1e8;
assign q[7623]= 16'hddd3;
assign q[7624]= 16'hd9db;
assign q[7625]= 16'hd613;
assign q[7626]= 16'hd28a;
assign q[7627]= 16'hcf52;
assign q[7628]= 16'hcc7a;
assign q[7629]= 16'hca0f;
assign q[7630]= 16'hc821;
assign q[7631]= 16'hc6b8;
assign q[7632]= 16'hc5df;
assign q[7633]= 16'hc59d;
assign q[7634]= 16'hc5f6;
assign q[7635]= 16'hc6eb;
assign q[7636]= 16'hc87a;
assign q[7637]= 16'hcaa0;
assign q[7638]= 16'hcd54;
assign q[7639]= 16'hd08c;
assign q[7640]= 16'hd439;
assign q[7641]= 16'hd84c;
assign q[7642]= 16'hdcb0;
assign q[7643]= 16'he150;
assign q[7644]= 16'he616;
assign q[7645]= 16'heae7;
assign q[7646]= 16'hefab;
assign q[7647]= 16'hf447;
assign q[7648]= 16'hf8a3;
assign q[7649]= 16'hfca6;
assign q[7650]= 16'h39;
assign q[7651]= 16'h348;
assign q[7652]= 16'h5c3;
assign q[7653]= 16'h79b;
assign q[7654]= 16'h8c6;
assign q[7655]= 16'h93f;
assign q[7656]= 16'h903;
assign q[7657]= 16'h817;
assign q[7658]= 16'h682;
assign q[7659]= 16'h450;
assign q[7660]= 16'h193;
assign q[7661]= 16'hfe5f;
assign q[7662]= 16'hfaca;
assign q[7663]= 16'hf6f0;
assign q[7664]= 16'hf2ec;
assign q[7665]= 16'heedb;
assign q[7666]= 16'headc;
assign q[7667]= 16'he70b;
assign q[7668]= 16'he384;
assign q[7669]= 16'he061;
assign q[7670]= 16'hddba;
assign q[7671]= 16'hdba1;
assign q[7672]= 16'hda27;
assign q[7673]= 16'hd956;
assign q[7674]= 16'hd937;
assign q[7675]= 16'hd9cb;
assign q[7676]= 16'hdb10;
assign q[7677]= 16'hdd00;
assign q[7678]= 16'hdf90;
assign q[7679]= 16'he2b2;
assign q[7680]= 16'he654;
assign q[7681]= 16'hea62;
assign q[7682]= 16'heec8;
assign q[7683]= 16'hf36d;
assign q[7684]= 16'hf83c;
assign q[7685]= 16'hfd1d;
assign q[7686]= 16'h1f9;
assign q[7687]= 16'h6bf;
assign q[7688]= 16'hb59;
assign q[7689]= 16'hfb9;
assign q[7690]= 16'h13d1;
assign q[7691]= 16'h1797;
assign q[7692]= 16'h1b02;
assign q[7693]= 16'h1e0e;
assign q[7694]= 16'h20b9;
assign q[7695]= 16'h2304;
assign q[7696]= 16'h24f2;
assign q[7697]= 16'h2687;
assign q[7698]= 16'h27c9;
assign q[7699]= 16'h28c1;
assign q[7700]= 16'h2977;
assign q[7701]= 16'h29f4;
assign q[7702]= 16'h2a40;
assign q[7703]= 16'h2a65;
assign q[7704]= 16'h2a6c;
assign q[7705]= 16'h2a5d;
assign q[7706]= 16'h2a3f;
assign q[7707]= 16'h2a19;
assign q[7708]= 16'h29f2;
assign q[7709]= 16'h29cd;
assign q[7710]= 16'h29b1;
assign q[7711]= 16'h29a1;
assign q[7712]= 16'h299f;
assign q[7713]= 16'h29af;
assign q[7714]= 16'h29d3;
assign q[7715]= 16'h2a0b;
assign q[7716]= 16'h2a59;
assign q[7717]= 16'h2abd;
assign q[7718]= 16'h2b36;
assign q[7719]= 16'h2bc3;
assign q[7720]= 16'h2c61;
assign q[7721]= 16'h2d0e;
assign q[7722]= 16'h2dc4;
assign q[7723]= 16'h2e80;
assign q[7724]= 16'h2f3a;
assign q[7725]= 16'h2feb;
assign q[7726]= 16'h308b;
assign q[7727]= 16'h3111;
assign q[7728]= 16'h3173;
assign q[7729]= 16'h31a6;
assign q[7730]= 16'h31a0;
assign q[7731]= 16'h3159;
assign q[7732]= 16'h30c5;
assign q[7733]= 16'h2fdd;
assign q[7734]= 16'h2e9b;
assign q[7735]= 16'h2cfa;
assign q[7736]= 16'h2af7;
assign q[7737]= 16'h2893;
assign q[7738]= 16'h25d0;
assign q[7739]= 16'h22b3;
assign q[7740]= 16'h1f47;
assign q[7741]= 16'h1b95;
assign q[7742]= 16'h17ac;
assign q[7743]= 16'h139c;
assign q[7744]= 16'hf77;
assign q[7745]= 16'hb50;
assign q[7746]= 16'h73b;
assign q[7747]= 16'h34a;
assign q[7748]= 16'hff93;
assign q[7749]= 16'hfc24;
assign q[7750]= 16'hf90d;
assign q[7751]= 16'hf65b;
assign q[7752]= 16'hf415;
assign q[7753]= 16'hf242;
assign q[7754]= 16'hf0e2;
assign q[7755]= 16'heff3;
assign q[7756]= 16'hef6c;
assign q[7757]= 16'hef44;
assign q[7758]= 16'hef6c;
assign q[7759]= 16'hefd2;
assign q[7760]= 16'hf063;
assign q[7761]= 16'hf10a;
assign q[7762]= 16'hf1b2;
assign q[7763]= 16'hf244;
assign q[7764]= 16'hf2ae;
assign q[7765]= 16'hf2dc;
assign q[7766]= 16'hf2c0;
assign q[7767]= 16'hf24e;
assign q[7768]= 16'hf17e;
assign q[7769]= 16'hf04f;
assign q[7770]= 16'heec1;
assign q[7771]= 16'hecdb;
assign q[7772]= 16'heaa9;
assign q[7773]= 16'he839;
assign q[7774]= 16'he59f;
assign q[7775]= 16'he2f0;
assign q[7776]= 16'he045;
assign q[7777]= 16'hddb6;
assign q[7778]= 16'hdb5d;
assign q[7779]= 16'hd953;
assign q[7780]= 16'hd7ad;
assign q[7781]= 16'hd680;
assign q[7782]= 16'hd5dd;
assign q[7783]= 16'hd5cf;
assign q[7784]= 16'hd65d;
assign q[7785]= 16'hd78c;
assign q[7786]= 16'hd956;
assign q[7787]= 16'hdbb6;
assign q[7788]= 16'hde9d;
assign q[7789]= 16'he1fb;
assign q[7790]= 16'he5bb;
assign q[7791]= 16'he9c6;
assign q[7792]= 16'hee00;
assign q[7793]= 16'hf24e;
assign q[7794]= 16'hf695;
assign q[7795]= 16'hfaba;
assign q[7796]= 16'hfea2;
assign q[7797]= 16'h235;
assign q[7798]= 16'h561;
assign q[7799]= 16'h814;
assign q[7800]= 16'ha41;
assign q[7801]= 16'hbdf;
assign q[7802]= 16'hcea;
assign q[7803]= 16'hd62;
assign q[7804]= 16'hd4a;
assign q[7805]= 16'hcaa;
assign q[7806]= 16'hb8e;
assign q[7807]= 16'ha03;
assign q[7808]= 16'h818;
assign q[7809]= 16'h5de;
assign q[7810]= 16'h369;
assign q[7811]= 16'hca;
assign q[7812]= 16'hfe15;
assign q[7813]= 16'hfb58;
assign q[7814]= 16'hf8a5;
assign q[7815]= 16'hf60b;
assign q[7816]= 16'hf396;
assign q[7817]= 16'hf153;
assign q[7818]= 16'hef4a;
assign q[7819]= 16'hed83;
assign q[7820]= 16'hec03;
assign q[7821]= 16'head0;
assign q[7822]= 16'he9eb;
assign q[7823]= 16'he956;
assign q[7824]= 16'he913;
assign q[7825]= 16'he920;
assign q[7826]= 16'he97c;
assign q[7827]= 16'hea26;
assign q[7828]= 16'heb19;
assign q[7829]= 16'hec54;
assign q[7830]= 16'hedd1;
assign q[7831]= 16'hef8c;
assign q[7832]= 16'hf17f;
assign q[7833]= 16'hf3a1;
assign q[7834]= 16'hf5ec;
assign q[7835]= 16'hf855;
assign q[7836]= 16'hfad3;
assign q[7837]= 16'hfd58;
assign q[7838]= 16'hffda;
assign q[7839]= 16'h249;
assign q[7840]= 16'h499;
assign q[7841]= 16'h6bb;
assign q[7842]= 16'h8a2;
assign q[7843]= 16'ha40;
assign q[7844]= 16'hb8a;
assign q[7845]= 16'hc74;
assign q[7846]= 16'hcf9;
assign q[7847]= 16'hd11;
assign q[7848]= 16'hcbc;
assign q[7849]= 16'hbfa;
assign q[7850]= 16'hacf;
assign q[7851]= 16'h945;
assign q[7852]= 16'h767;
assign q[7853]= 16'h544;
assign q[7854]= 16'h2f0;
assign q[7855]= 16'h7e;
assign q[7856]= 16'hfe06;
assign q[7857]= 16'hfb9f;
assign q[7858]= 16'hf961;
assign q[7859]= 16'hf765;
assign q[7860]= 16'hf5c0;
assign q[7861]= 16'hf488;
assign q[7862]= 16'hf3ce;
assign q[7863]= 16'hf3a0;
assign q[7864]= 16'hf407;
assign q[7865]= 16'hf508;
assign q[7866]= 16'hf6a4;
assign q[7867]= 16'hf8d6;
assign q[7868]= 16'hfb93;
assign q[7869]= 16'hfecf;
assign q[7870]= 16'h276;
assign q[7871]= 16'h675;
assign q[7872]= 16'hab1;
assign q[7873]= 16'hf13;
assign q[7874]= 16'h137e;
assign q[7875]= 16'h17d9;
assign q[7876]= 16'h1c0b;
assign q[7877]= 16'h1ffc;
assign q[7878]= 16'h2398;
assign q[7879]= 16'h26ce;
assign q[7880]= 16'h2993;
assign q[7881]= 16'h2bde;
assign q[7882]= 16'h2dab;
assign q[7883]= 16'h2efd;
assign q[7884]= 16'h2fd8;
assign q[7885]= 16'h3047;
assign q[7886]= 16'h3057;
assign q[7887]= 16'h3018;
assign q[7888]= 16'h2f9c;
assign q[7889]= 16'h2ef6;
assign q[7890]= 16'h2e3a;
assign q[7891]= 16'h2d7a;
assign q[7892]= 16'h2cc7;
assign q[7893]= 16'h2c31;
assign q[7894]= 16'h2bc4;
assign q[7895]= 16'h2b87;
assign q[7896]= 16'h2b80;
assign q[7897]= 16'h2baf;
assign q[7898]= 16'h2c12;
assign q[7899]= 16'h2ca1;
assign q[7900]= 16'h2d52;
assign q[7901]= 16'h2e18;
assign q[7902]= 16'h2ee3;
assign q[7903]= 16'h2fa2;
assign q[7904]= 16'h3042;
assign q[7905]= 16'h30b1;
assign q[7906]= 16'h30de;
assign q[7907]= 16'h30b7;
assign q[7908]= 16'h302d;
assign q[7909]= 16'h2f35;
assign q[7910]= 16'h2dc5;
assign q[7911]= 16'h2bd6;
assign q[7912]= 16'h2966;
assign q[7913]= 16'h2674;
assign q[7914]= 16'h2305;
assign q[7915]= 16'h1f1e;
assign q[7916]= 16'h1acb;
assign q[7917]= 16'h1616;
assign q[7918]= 16'h110d;
assign q[7919]= 16'hbc1;
assign q[7920]= 16'h641;
assign q[7921]= 16'h9e;
assign q[7922]= 16'hfaec;
assign q[7923]= 16'hf53a;
assign q[7924]= 16'hef99;
assign q[7925]= 16'hea1a;
assign q[7926]= 16'he4cc;
assign q[7927]= 16'hdfbe;
assign q[7928]= 16'hdafe;
assign q[7929]= 16'hd697;
assign q[7930]= 16'hd296;
assign q[7931]= 16'hcf06;
assign q[7932]= 16'hcbef;
assign q[7933]= 16'hc95b;
assign q[7934]= 16'hc751;
assign q[7935]= 16'hc5d7;
assign q[7936]= 16'hc4f4;
assign q[7937]= 16'hc4ac;
assign q[7938]= 16'hc501;
assign q[7939]= 16'hc5f3;
assign q[7940]= 16'hc782;
assign q[7941]= 16'hc9aa;
assign q[7942]= 16'hcc65;
assign q[7943]= 16'hcfa9;
assign q[7944]= 16'hd36a;
assign q[7945]= 16'hd79a;
assign q[7946]= 16'hdc26;
assign q[7947]= 16'he0f9;
assign q[7948]= 16'he5fb;
assign q[7949]= 16'heb12;
assign q[7950]= 16'hf023;
assign q[7951]= 16'hf510;
assign q[7952]= 16'hf9bd;
assign q[7953]= 16'hfe0b;
assign q[7954]= 16'h1df;
assign q[7955]= 16'h522;
assign q[7956]= 16'h7bd;
assign q[7957]= 16'h99c;
assign q[7958]= 16'hab5;
assign q[7959]= 16'hafd;
assign q[7960]= 16'ha75;
assign q[7961]= 16'h91f;
assign q[7962]= 16'h707;
assign q[7963]= 16'h43e;
assign q[7964]= 16'hda;
assign q[7965]= 16'hfcf7;
assign q[7966]= 16'hf8b5;
assign q[7967]= 16'hf437;
assign q[7968]= 16'hefa4;
assign q[7969]= 16'heb23;
assign q[7970]= 16'he6d9;
assign q[7971]= 16'he2ed;
assign q[7972]= 16'hdf80;
assign q[7973]= 16'hdcaf;
assign q[7974]= 16'hda94;
assign q[7975]= 16'hd942;
assign q[7976]= 16'hd8c2;
assign q[7977]= 16'hd91b;
assign q[7978]= 16'hda48;
assign q[7979]= 16'hdc3f;
assign q[7980]= 16'hdeef;
assign q[7981]= 16'he23f;
assign q[7982]= 16'he612;
assign q[7983]= 16'hea46;
assign q[7984]= 16'heeb5;
assign q[7985]= 16'hf338;
assign q[7986]= 16'hf7a7;
assign q[7987]= 16'hfbdc;
assign q[7988]= 16'hffb2;
assign q[7989]= 16'h306;
assign q[7990]= 16'h5bf;
assign q[7991]= 16'h7c4;
assign q[7992]= 16'h905;
assign q[7993]= 16'h978;
assign q[7994]= 16'h91b;
assign q[7995]= 16'h7f1;
assign q[7996]= 16'h606;
assign q[7997]= 16'h36b;
assign q[7998]= 16'h37;
assign q[7999]= 16'hfc85;
assign q[8000]= 16'hf873;
assign q[8001]= 16'hf424;
assign q[8002]= 16'hefba;
assign q[8003]= 16'heb58;
assign q[8004]= 16'he721;
assign q[8005]= 16'he335;
assign q[8006]= 16'hdfb1;
assign q[8007]= 16'hdcb1;
assign q[8008]= 16'hda4a;
assign q[8009]= 16'hd88d;
assign q[8010]= 16'hd788;
assign q[8011]= 16'hd743;
assign q[8012]= 16'hd7c2;
assign q[8013]= 16'hd902;
assign q[8014]= 16'hdaff;
assign q[8015]= 16'hddb0;
assign q[8016]= 16'he108;
assign q[8017]= 16'he4f7;
assign q[8018]= 16'he96c;
assign q[8019]= 16'hee53;
assign q[8020]= 16'hf396;
assign q[8021]= 16'hf921;
assign q[8022]= 16'hfedb;
assign q[8023]= 16'h4ad;
assign q[8024]= 16'ha82;
assign q[8025]= 16'h1040;
assign q[8026]= 16'h15d2;
assign q[8027]= 16'h1b21;
assign q[8028]= 16'h2017;
assign q[8029]= 16'h249e;
assign q[8030]= 16'h28a3;
assign q[8031]= 16'h2c12;
assign q[8032]= 16'h2edb;
assign q[8033]= 16'h30ee;
assign q[8034]= 16'h323d;
assign q[8035]= 16'h32be;
assign q[8036]= 16'h326a;
assign q[8037]= 16'h313c;
assign q[8038]= 16'h2f35;
assign q[8039]= 16'h2c5a;
assign q[8040]= 16'h28b3;
assign q[8041]= 16'h244e;
assign q[8042]= 16'h1f3f;
assign q[8043]= 16'h199e;
assign q[8044]= 16'h1387;
assign q[8045]= 16'hd1b;
assign q[8046]= 16'h67f;
assign q[8047]= 16'hffdb;
assign q[8048]= 16'hf956;
assign q[8049]= 16'hf31b;
assign q[8050]= 16'hed54;
assign q[8051]= 16'he827;
assign q[8052]= 16'he3bb;
assign q[8053]= 16'he02f;
assign q[8054]= 16'hdd9f;
assign q[8055]= 16'hdc1f;
assign q[8056]= 16'hdbbb;
assign q[8057]= 16'hdc7a;
assign q[8058]= 16'hde56;
assign q[8059]= 16'he143;
assign q[8060]= 16'he52c;
assign q[8061]= 16'he9f3;
assign q[8062]= 16'hef75;
assign q[8063]= 16'hf584;
assign q[8064]= 16'hfbf2;
assign q[8065]= 16'h289;
assign q[8066]= 16'h916;
assign q[8067]= 16'hf62;
assign q[8068]= 16'h1538;
assign q[8069]= 16'h1a67;
assign q[8070]= 16'h1ec4;
assign q[8071]= 16'h2228;
assign q[8072]= 16'h2477;
assign q[8073]= 16'h259b;
assign q[8074]= 16'h2588;
assign q[8075]= 16'h243e;
assign q[8076]= 16'h21c3;
assign q[8077]= 16'h1e2a;
assign q[8078]= 16'h198c;
assign q[8079]= 16'h140b;
assign q[8080]= 16'hdd0;
assign q[8081]= 16'h708;
assign q[8082]= 16'hffe3;
assign q[8083]= 16'hf891;
assign q[8084]= 16'hf145;
assign q[8085]= 16'hea2e;
assign q[8086]= 16'he378;
assign q[8087]= 16'hdd49;
assign q[8088]= 16'hd7c2;
assign q[8089]= 16'hd2fb;
assign q[8090]= 16'hcf07;
assign q[8091]= 16'hcbef;
assign q[8092]= 16'hc9b4;
assign q[8093]= 16'hc84f;
assign q[8094]= 16'hc7b5;
assign q[8095]= 16'hc7d0;
assign q[8096]= 16'hc889;
assign q[8097]= 16'hc9c5;
assign q[8098]= 16'hcb66;
assign q[8099]= 16'hcd4d;
assign q[8100]= 16'hcf5c;
assign q[8101]= 16'hd178;
assign q[8102]= 16'hd388;
assign q[8103]= 16'hd578;
assign q[8104]= 16'hd739;
assign q[8105]= 16'hd8c2;
assign q[8106]= 16'hda0d;
assign q[8107]= 16'hdb1e;
assign q[8108]= 16'hdbfb;
assign q[8109]= 16'hdcb0;
assign q[8110]= 16'hdd4e;
assign q[8111]= 16'hdde7;
assign q[8112]= 16'hde90;
assign q[8113]= 16'hdf5e;
assign q[8114]= 16'he068;
assign q[8115]= 16'he1c1;
assign q[8116]= 16'he379;
assign q[8117]= 16'he59d;
assign q[8118]= 16'he837;
assign q[8119]= 16'heb4a;
assign q[8120]= 16'heed5;
assign q[8121]= 16'hf2cf;
assign q[8122]= 16'hf72d;
assign q[8123]= 16'hfbdc;
assign q[8124]= 16'hc7;
assign q[8125]= 16'h5d3;
assign q[8126]= 16'hae5;
assign q[8127]= 16'hfde;
assign q[8128]= 16'h149e;
assign q[8129]= 16'h1906;
assign q[8130]= 16'h1cf9;
assign q[8131]= 16'h205c;
assign q[8132]= 16'h2317;
assign q[8133]= 16'h2517;
assign q[8134]= 16'h264b;
assign q[8135]= 16'h26ac;
assign q[8136]= 16'h2633;
assign q[8137]= 16'h24e2;
assign q[8138]= 16'h22bf;
assign q[8139]= 16'h1fd5;
assign q[8140]= 16'h1c33;
assign q[8141]= 16'h17ec;
assign q[8142]= 16'h1317;
assign q[8143]= 16'hdcd;
assign q[8144]= 16'h829;
assign q[8145]= 16'h246;
assign q[8146]= 16'hfc40;
assign q[8147]= 16'hf632;
assign q[8148]= 16'hf037;
assign q[8149]= 16'hea65;
assign q[8150]= 16'he4d5;
assign q[8151]= 16'hdf9a;
assign q[8152]= 16'hdac5;
assign q[8153]= 16'hd664;
assign q[8154]= 16'hd283;
assign q[8155]= 16'hcf2b;
assign q[8156]= 16'hcc61;
assign q[8157]= 16'hca2a;
assign q[8158]= 16'hc885;
assign q[8159]= 16'hc772;
assign q[8160]= 16'hc6ed;
assign q[8161]= 16'hc6f1;
assign q[8162]= 16'hc778;
assign q[8163]= 16'hc879;
assign q[8164]= 16'hc9eb;
assign q[8165]= 16'hcbc1;
assign q[8166]= 16'hcdf1;
assign q[8167]= 16'hd06d;
assign q[8168]= 16'hd327;
assign q[8169]= 16'hd610;
assign q[8170]= 16'hd918;
assign q[8171]= 16'hdc2e;
assign q[8172]= 16'hdf43;
assign q[8173]= 16'he244;
assign q[8174]= 16'he523;
assign q[8175]= 16'he7cd;
assign q[8176]= 16'hea33;
assign q[8177]= 16'hec49;
assign q[8178]= 16'hee00;
assign q[8179]= 16'hef4d;
assign q[8180]= 16'hf02a;
assign q[8181]= 16'hf090;
assign q[8182]= 16'hf07d;
assign q[8183]= 16'heff2;
assign q[8184]= 16'heef3;
assign q[8185]= 16'hed89;
assign q[8186]= 16'hebbe;
assign q[8187]= 16'he9a2;
assign q[8188]= 16'he747;
assign q[8189]= 16'he4c1;
assign q[8190]= 16'he228;
assign q[8191]= 16'hdf93;
assign q[8192]= 16'hdd1d;
assign q[8193]= 16'hdae0;
assign q[8194]= 16'hd8f4;
assign q[8195]= 16'hd771;
assign q[8196]= 16'hd66d;
assign q[8197]= 16'hd5fb;
assign q[8198]= 16'hd62a;
assign q[8199]= 16'hd705;
assign q[8200]= 16'hd894;
assign q[8201]= 16'hdad8;
assign q[8202]= 16'hddce;
assign q[8203]= 16'he16e;
assign q[8204]= 16'he5ab;
assign q[8205]= 16'hea74;
assign q[8206]= 16'hefb3;
assign q[8207]= 16'hf54f;
assign q[8208]= 16'hfb2c;
assign q[8209]= 16'h12d;
assign q[8210]= 16'h732;
assign q[8211]= 16'hd1d;
assign q[8212]= 16'h12cf;
assign q[8213]= 16'h182b;
assign q[8214]= 16'h1d16;
assign q[8215]= 16'h2178;
assign q[8216]= 16'h253e;
assign q[8217]= 16'h2857;
assign q[8218]= 16'h2ab9;
assign q[8219]= 16'h2c5e;
assign q[8220]= 16'h2d43;
assign q[8221]= 16'h2d6b;
assign q[8222]= 16'h2cdf;
assign q[8223]= 16'h2baa;
assign q[8224]= 16'h29db;
assign q[8225]= 16'h2786;
assign q[8226]= 16'h24bd;
assign q[8227]= 16'h2199;
assign q[8228]= 16'h1e2f;
assign q[8229]= 16'h1a97;
assign q[8230]= 16'h16e9;
assign q[8231]= 16'h1338;
assign q[8232]= 16'hf9a;
assign q[8233]= 16'hc1e;
assign q[8234]= 16'h8d4;
assign q[8235]= 16'h5c6;
assign q[8236]= 16'h2fe;
assign q[8237]= 16'h80;
assign q[8238]= 16'hfe50;
assign q[8239]= 16'hfc6a;
assign q[8240]= 16'hfacd;
assign q[8241]= 16'hf973;
assign q[8242]= 16'hf854;
assign q[8243]= 16'hf768;
assign q[8244]= 16'hf6a7;
assign q[8245]= 16'hf605;
assign q[8246]= 16'hf57b;
assign q[8247]= 16'hf4ff;
assign q[8248]= 16'hf48b;
assign q[8249]= 16'hf418;
assign q[8250]= 16'hf3a2;
assign q[8251]= 16'hf325;
assign q[8252]= 16'hf2a2;
assign q[8253]= 16'hf219;
assign q[8254]= 16'hf18b;
assign q[8255]= 16'hf0fe;
assign q[8256]= 16'hf075;
assign q[8257]= 16'heff6;
assign q[8258]= 16'hef87;
assign q[8259]= 16'hef2d;
assign q[8260]= 16'heeed;
assign q[8261]= 16'heecc;
assign q[8262]= 16'heecc;
assign q[8263]= 16'heef0;
assign q[8264]= 16'hef38;
assign q[8265]= 16'hefa1;
assign q[8266]= 16'hf028;
assign q[8267]= 16'hf0c8;
assign q[8268]= 16'hf179;
assign q[8269]= 16'hf234;
assign q[8270]= 16'hf2f0;
assign q[8271]= 16'hf3a1;
assign q[8272]= 16'hf440;
assign q[8273]= 16'hf4c1;
assign q[8274]= 16'hf51c;
assign q[8275]= 16'hf549;
assign q[8276]= 16'hf543;
assign q[8277]= 16'hf505;
assign q[8278]= 16'hf48e;
assign q[8279]= 16'hf3e0;
assign q[8280]= 16'hf2fd;
assign q[8281]= 16'hf1ef;
assign q[8282]= 16'hf0bc;
assign q[8283]= 16'hef73;
assign q[8284]= 16'hee21;
assign q[8285]= 16'hecd5;
assign q[8286]= 16'heba2;
assign q[8287]= 16'hea99;
assign q[8288]= 16'he9cc;
assign q[8289]= 16'he94b;
assign q[8290]= 16'he926;
assign q[8291]= 16'he96c;
assign q[8292]= 16'hea27;
assign q[8293]= 16'heb5e;
assign q[8294]= 16'hed17;
assign q[8295]= 16'hef51;
assign q[8296]= 16'hf208;
assign q[8297]= 16'hf535;
assign q[8298]= 16'hf8cb;
assign q[8299]= 16'hfcbb;
assign q[8300]= 16'hf1;
assign q[8301]= 16'h558;
assign q[8302]= 16'h9d7;
assign q[8303]= 16'he54;
assign q[8304]= 16'h12b4;
assign q[8305]= 16'h16dc;
assign q[8306]= 16'h1ab4;
assign q[8307]= 16'h1e21;
assign q[8308]= 16'h2110;
assign q[8309]= 16'h236d;
assign q[8310]= 16'h2529;
assign q[8311]= 16'h263a;
assign q[8312]= 16'h269a;
assign q[8313]= 16'h2648;
assign q[8314]= 16'h2546;
assign q[8315]= 16'h239e;
assign q[8316]= 16'h215c;
assign q[8317]= 16'h1e90;
assign q[8318]= 16'h1b4e;
assign q[8319]= 16'h17ad;
assign q[8320]= 16'h13c6;
assign q[8321]= 16'hfb4;
assign q[8322]= 16'hb91;
assign q[8323]= 16'h779;
assign q[8324]= 16'h385;
assign q[8325]= 16'hffce;
assign q[8326]= 16'hfc69;
assign q[8327]= 16'hf969;
assign q[8328]= 16'hf6e0;
assign q[8329]= 16'hf4d8;
assign q[8330]= 16'hf35b;
assign q[8331]= 16'hf26e;
assign q[8332]= 16'hf213;
assign q[8333]= 16'hf245;
assign q[8334]= 16'hf300;
assign q[8335]= 16'hf43b;
assign q[8336]= 16'hf5e9;
assign q[8337]= 16'hf7fd;
assign q[8338]= 16'hfa68;
assign q[8339]= 16'hfd17;
assign q[8340]= 16'hfff9;
assign q[8341]= 16'h2fa;
assign q[8342]= 16'h60a;
assign q[8343]= 16'h917;
assign q[8344]= 16'hc0d;
assign q[8345]= 16'hedd;
assign q[8346]= 16'h1178;
assign q[8347]= 16'h13cf;
assign q[8348]= 16'h15d7;
assign q[8349]= 16'h1784;
assign q[8350]= 16'h18cc;
assign q[8351]= 16'h19a9;
assign q[8352]= 16'h1a15;
assign q[8353]= 16'h1a0c;
assign q[8354]= 16'h198a;
assign q[8355]= 16'h1891;
assign q[8356]= 16'h1721;
assign q[8357]= 16'h153d;
assign q[8358]= 16'h12eb;
assign q[8359]= 16'h1031;
assign q[8360]= 16'hd18;
assign q[8361]= 16'h9ab;
assign q[8362]= 16'h5f5;
assign q[8363]= 16'h205;
assign q[8364]= 16'hfdeb;
assign q[8365]= 16'hf9b6;
assign q[8366]= 16'hf57a;
assign q[8367]= 16'hf149;
assign q[8368]= 16'hed37;
assign q[8369]= 16'he957;
assign q[8370]= 16'he5bd;
assign q[8371]= 16'he27c;
assign q[8372]= 16'hdfa5;
assign q[8373]= 16'hdd48;
assign q[8374]= 16'hdb73;
assign q[8375]= 16'hda31;
assign q[8376]= 16'hd98a;
assign q[8377]= 16'hd983;
assign q[8378]= 16'hda1e;
assign q[8379]= 16'hdb59;
assign q[8380]= 16'hdd2f;
assign q[8381]= 16'hdf96;
assign q[8382]= 16'he282;
assign q[8383]= 16'he5e4;
assign q[8384]= 16'he9aa;
assign q[8385]= 16'hedc0;
assign q[8386]= 16'hf211;
assign q[8387]= 16'hf687;
assign q[8388]= 16'hfb0d;
assign q[8389]= 16'hff8d;
assign q[8390]= 16'h3f2;
assign q[8391]= 16'h82b;
assign q[8392]= 16'hc2a;
assign q[8393]= 16'hfe0;
assign q[8394]= 16'h1345;
assign q[8395]= 16'h1653;
assign q[8396]= 16'h1908;
assign q[8397]= 16'h1b65;
assign q[8398]= 16'h1d6f;
assign q[8399]= 16'h1f2e;
assign q[8400]= 16'h20aa;
assign q[8401]= 16'h21f1;
assign q[8402]= 16'h230f;
assign q[8403]= 16'h2411;
assign q[8404]= 16'h2505;
assign q[8405]= 16'h25f6;
assign q[8406]= 16'h26ef;
assign q[8407]= 16'h27f8;
assign q[8408]= 16'h2916;
assign q[8409]= 16'h2a4b;
assign q[8410]= 16'h2b96;
assign q[8411]= 16'h2cf1;
assign q[8412]= 16'h2e54;
assign q[8413]= 16'h2fb4;
assign q[8414]= 16'h3101;
assign q[8415]= 16'h322c;
assign q[8416]= 16'h3321;
assign q[8417]= 16'h33ce;
assign q[8418]= 16'h3420;
assign q[8419]= 16'h3404;
assign q[8420]= 16'h3369;
assign q[8421]= 16'h3242;
assign q[8422]= 16'h3083;
assign q[8423]= 16'h2e26;
assign q[8424]= 16'h2b27;
assign q[8425]= 16'h278a;
assign q[8426]= 16'h2353;
assign q[8427]= 16'h1e90;
assign q[8428]= 16'h1951;
assign q[8429]= 16'h13a9;
assign q[8430]= 16'hdb1;
assign q[8431]= 16'h784;
assign q[8432]= 16'h13f;
assign q[8433]= 16'hfb02;
assign q[8434]= 16'hf4e9;
assign q[8435]= 16'hef13;
assign q[8436]= 16'he99e;
assign q[8437]= 16'he4a2;
assign q[8438]= 16'he037;
assign q[8439]= 16'hdc6e;
assign q[8440]= 16'hd957;
assign q[8441]= 16'hd6f9;
assign q[8442]= 16'hd55a;
assign q[8443]= 16'hd478;
assign q[8444]= 16'hd44c;
assign q[8445]= 16'hd4cd;
assign q[8446]= 16'hd5ec;
assign q[8447]= 16'hd797;
assign q[8448]= 16'hd9b9;
assign q[8449]= 16'hdc3b;
assign q[8450]= 16'hdf06;
assign q[8451]= 16'he203;
assign q[8452]= 16'he51b;
assign q[8453]= 16'he839;
assign q[8454]= 16'heb4a;
assign q[8455]= 16'hee3d;
assign q[8456]= 16'hf107;
assign q[8457]= 16'hf39d;
assign q[8458]= 16'hf5fb;
assign q[8459]= 16'hf81e;
assign q[8460]= 16'hfa0a;
assign q[8461]= 16'hfbc2;
assign q[8462]= 16'hfd4e;
assign q[8463]= 16'hfeb8;
assign q[8464]= 16'hb;
assign q[8465]= 16'h155;
assign q[8466]= 16'h2a2;
assign q[8467]= 16'h3fd;
assign q[8468]= 16'h572;
assign q[8469]= 16'h709;
assign q[8470]= 16'h8c9;
assign q[8471]= 16'hab7;
assign q[8472]= 16'hcd3;
assign q[8473]= 16'hf1d;
assign q[8474]= 16'h118e;
assign q[8475]= 16'h1420;
assign q[8476]= 16'h16c9;
assign q[8477]= 16'h197b;
assign q[8478]= 16'h1c28;
assign q[8479]= 16'h1ec0;
assign q[8480]= 16'h2134;
assign q[8481]= 16'h2373;
assign q[8482]= 16'h256c;
assign q[8483]= 16'h2711;
assign q[8484]= 16'h2854;
assign q[8485]= 16'h292a;
assign q[8486]= 16'h298a;
assign q[8487]= 16'h296e;
assign q[8488]= 16'h28d3;
assign q[8489]= 16'h27b7;
assign q[8490]= 16'h261f;
assign q[8491]= 16'h2410;
assign q[8492]= 16'h2191;
assign q[8493]= 16'h1eae;
assign q[8494]= 16'h1b73;
assign q[8495]= 16'h17ee;
assign q[8496]= 16'h1430;
assign q[8497]= 16'h1048;
assign q[8498]= 16'hc47;
assign q[8499]= 16'h83e;
assign q[8500]= 16'h43e;
assign q[8501]= 16'h56;
assign q[8502]= 16'hfc95;
assign q[8503]= 16'hf908;
assign q[8504]= 16'hf5ba;
assign q[8505]= 16'hf2b7;
assign q[8506]= 16'hf008;
assign q[8507]= 16'hedb3;
assign q[8508]= 16'hebbe;
assign q[8509]= 16'hea2c;
assign q[8510]= 16'he901;
assign q[8511]= 16'he83e;
assign q[8512]= 16'he7e0;
assign q[8513]= 16'he7e8;
assign q[8514]= 16'he851;
assign q[8515]= 16'he918;
assign q[8516]= 16'hea36;
assign q[8517]= 16'heba6;
assign q[8518]= 16'hed61;
assign q[8519]= 16'hef5c;
assign q[8520]= 16'hf18f;
assign q[8521]= 16'hf3f0;
assign q[8522]= 16'hf672;
assign q[8523]= 16'hf90a;
assign q[8524]= 16'hfbab;
assign q[8525]= 16'hfe46;
assign q[8526]= 16'hce;
assign q[8527]= 16'h336;
assign q[8528]= 16'h56f;
assign q[8529]= 16'h76b;
assign q[8530]= 16'h91d;
assign q[8531]= 16'ha79;
assign q[8532]= 16'hb74;
assign q[8533]= 16'hc05;
assign q[8534]= 16'hc25;
assign q[8535]= 16'hbce;
assign q[8536]= 16'hafd;
assign q[8537]= 16'h9b2;
assign q[8538]= 16'h7ef;
assign q[8539]= 16'h5ba;
assign q[8540]= 16'h31a;
assign q[8541]= 16'h18;
assign q[8542]= 16'hfcc4;
assign q[8543]= 16'hf929;
assign q[8544]= 16'hf558;
assign q[8545]= 16'hf162;
assign q[8546]= 16'hed5b;
assign q[8547]= 16'he953;
assign q[8548]= 16'he55f;
assign q[8549]= 16'he18e;
assign q[8550]= 16'hddf1;
assign q[8551]= 16'hda98;
assign q[8552]= 16'hd78e;
assign q[8553]= 16'hd4de;
assign q[8554]= 16'hd28f;
assign q[8555]= 16'hd0a6;
assign q[8556]= 16'hcf27;
assign q[8557]= 16'hce0f;
assign q[8558]= 16'hcd5d;
assign q[8559]= 16'hcd0b;
assign q[8560]= 16'hcd12;
assign q[8561]= 16'hcd69;
assign q[8562]= 16'hce06;
assign q[8563]= 16'hcedf;
assign q[8564]= 16'hcfe8;
assign q[8565]= 16'hd118;
assign q[8566]= 16'hd263;
assign q[8567]= 16'hd3c1;
assign q[8568]= 16'hd52a;
assign q[8569]= 16'hd698;
assign q[8570]= 16'hd807;
assign q[8571]= 16'hd974;
assign q[8572]= 16'hdadf;
assign q[8573]= 16'hdc47;
assign q[8574]= 16'hddaf;
assign q[8575]= 16'hdf1b;
assign q[8576]= 16'he08f;
assign q[8577]= 16'he210;
assign q[8578]= 16'he3a2;
assign q[8579]= 16'he54b;
assign q[8580]= 16'he70e;
assign q[8581]= 16'he8ef;
assign q[8582]= 16'heaf0;
assign q[8583]= 16'hed11;
assign q[8584]= 16'hef50;
assign q[8585]= 16'hf1ab;
assign q[8586]= 16'hf41d;
assign q[8587]= 16'hf69f;
assign q[8588]= 16'hf92a;
assign q[8589]= 16'hfbb4;
assign q[8590]= 16'hfe33;
assign q[8591]= 16'h9c;
assign q[8592]= 16'h2e5;
assign q[8593]= 16'h503;
assign q[8594]= 16'h6ec;
assign q[8595]= 16'h896;
assign q[8596]= 16'h9f8;
assign q[8597]= 16'hb0d;
assign q[8598]= 16'hbcf;
assign q[8599]= 16'hc3c;
assign q[8600]= 16'hc52;
assign q[8601]= 16'hc13;
assign q[8602]= 16'hb82;
assign q[8603]= 16'haa4;
assign q[8604]= 16'h97f;
assign q[8605]= 16'h81c;
assign q[8606]= 16'h683;
assign q[8607]= 16'h4bf;
assign q[8608]= 16'h2da;
assign q[8609]= 16'hdf;
assign q[8610]= 16'hfed8;
assign q[8611]= 16'hfccf;
assign q[8612]= 16'hface;
assign q[8613]= 16'hf8dd;
assign q[8614]= 16'hf703;
assign q[8615]= 16'hf548;
assign q[8616]= 16'hf3b1;
assign q[8617]= 16'hf242;
assign q[8618]= 16'hf0fd;
assign q[8619]= 16'hefe5;
assign q[8620]= 16'heefc;
assign q[8621]= 16'hee40;
assign q[8622]= 16'hedb3;
assign q[8623]= 16'hed52;
assign q[8624]= 16'hed1c;
assign q[8625]= 16'hed10;
assign q[8626]= 16'hed2a;
assign q[8627]= 16'hed69;
assign q[8628]= 16'hedc9;
assign q[8629]= 16'hee47;
assign q[8630]= 16'heee0;
assign q[8631]= 16'hef90;
assign q[8632]= 16'hf051;
assign q[8633]= 16'hf120;
assign q[8634]= 16'hf1f6;
assign q[8635]= 16'hf2cd;
assign q[8636]= 16'hf39f;
assign q[8637]= 16'hf465;
assign q[8638]= 16'hf515;
assign q[8639]= 16'hf5aa;
assign q[8640]= 16'hf61a;
assign q[8641]= 16'hf65d;
assign q[8642]= 16'hf66d;
assign q[8643]= 16'hf642;
assign q[8644]= 16'hf5d7;
assign q[8645]= 16'hf526;
assign q[8646]= 16'hf42e;
assign q[8647]= 16'hf2ee;
assign q[8648]= 16'hf167;
assign q[8649]= 16'hef9c;
assign q[8650]= 16'hed95;
assign q[8651]= 16'heb58;
assign q[8652]= 16'he8f2;
assign q[8653]= 16'he670;
assign q[8654]= 16'he3e0;
assign q[8655]= 16'he152;
assign q[8656]= 16'hded8;
assign q[8657]= 16'hdc84;
assign q[8658]= 16'hda66;
assign q[8659]= 16'hd890;
assign q[8660]= 16'hd710;
assign q[8661]= 16'hd5f4;
assign q[8662]= 16'hd546;
assign q[8663]= 16'hd50b;
assign q[8664]= 16'hd549;
assign q[8665]= 16'hd5fd;
assign q[8666]= 16'hd722;
assign q[8667]= 16'hd8b1;
assign q[8668]= 16'hda9c;
assign q[8669]= 16'hdcd2;
assign q[8670]= 16'hdf3f;
assign q[8671]= 16'he1ce;
assign q[8672]= 16'he466;
assign q[8673]= 16'he6ee;
assign q[8674]= 16'he94d;
assign q[8675]= 16'heb6c;
assign q[8676]= 16'hed34;
assign q[8677]= 16'hee92;
assign q[8678]= 16'hef77;
assign q[8679]= 16'hefd7;
assign q[8680]= 16'hefad;
assign q[8681]= 16'heef8;
assign q[8682]= 16'hedbd;
assign q[8683]= 16'hec07;
assign q[8684]= 16'he9e5;
assign q[8685]= 16'he76d;
assign q[8686]= 16'he4b9;
assign q[8687]= 16'he1e6;
assign q[8688]= 16'hdf12;
assign q[8689]= 16'hdc61;
assign q[8690]= 16'hd9f2;
assign q[8691]= 16'hd7e7;
assign q[8692]= 16'hd65e;
assign q[8693]= 16'hd573;
assign q[8694]= 16'hd53b;
assign q[8695]= 16'hd5c9;
assign q[8696]= 16'hd727;
assign q[8697]= 16'hd95a;
assign q[8698]= 16'hdc61;
assign q[8699]= 16'he032;
assign q[8700]= 16'he4bd;
assign q[8701]= 16'he9ec;
assign q[8702]= 16'hefa2;
assign q[8703]= 16'hf5c0;
assign q[8704]= 16'hfc21;
assign q[8705]= 16'h29c;
assign q[8706]= 16'h90d;
assign q[8707]= 16'hf4b;
assign q[8708]= 16'h1530;
assign q[8709]= 16'h1a98;
assign q[8710]= 16'h1f66;
assign q[8711]= 16'h237f;
assign q[8712]= 16'h26cf;
assign q[8713]= 16'h294a;
assign q[8714]= 16'h2aeb;
assign q[8715]= 16'h2bb1;
assign q[8716]= 16'h2ba6;
assign q[8717]= 16'h2ad9;
assign q[8718]= 16'h295f;
assign q[8719]= 16'h2753;
assign q[8720]= 16'h24d2;
assign q[8721]= 16'h21fe;
assign q[8722]= 16'h1efa;
assign q[8723]= 16'h1bea;
assign q[8724]= 16'h18f0;
assign q[8725]= 16'h162d;
assign q[8726]= 16'h13bd;
assign q[8727]= 16'h11ba;
assign q[8728]= 16'h1037;
assign q[8729]= 16'hf42;
assign q[8730]= 16'hee4;
assign q[8731]= 16'hf1d;
assign q[8732]= 16'hfea;
assign q[8733]= 16'h1142;
assign q[8734]= 16'h1315;
assign q[8735]= 16'h1550;
assign q[8736]= 16'h17de;
assign q[8737]= 16'h1aa5;
assign q[8738]= 16'h1d8b;
assign q[8739]= 16'h2076;
assign q[8740]= 16'h234e;
assign q[8741]= 16'h25fc;
assign q[8742]= 16'h286b;
assign q[8743]= 16'h2a8a;
assign q[8744]= 16'h2c4e;
assign q[8745]= 16'h2daf;
assign q[8746]= 16'h2eaa;
assign q[8747]= 16'h2f40;
assign q[8748]= 16'h2f79;
assign q[8749]= 16'h2f5e;
assign q[8750]= 16'h2efc;
assign q[8751]= 16'h2e65;
assign q[8752]= 16'h2daa;
assign q[8753]= 16'h2cdd;
assign q[8754]= 16'h2c12;
assign q[8755]= 16'h2b5b;
assign q[8756]= 16'h2ac6;
assign q[8757]= 16'h2a61;
assign q[8758]= 16'h2a37;
assign q[8759]= 16'h2a4c;
assign q[8760]= 16'h2aa3;
assign q[8761]= 16'h2b39;
assign q[8762]= 16'h2c08;
assign q[8763]= 16'h2d05;
assign q[8764]= 16'h2e22;
assign q[8765]= 16'h2f4e;
assign q[8766]= 16'h3075;
assign q[8767]= 16'h3183;
assign q[8768]= 16'h3261;
assign q[8769]= 16'h32fa;
assign q[8770]= 16'h3339;
assign q[8771]= 16'h330d;
assign q[8772]= 16'h3264;
assign q[8773]= 16'h3132;
assign q[8774]= 16'h2f6f;
assign q[8775]= 16'h2d14;
assign q[8776]= 16'h2a21;
assign q[8777]= 16'h269b;
assign q[8778]= 16'h2289;
assign q[8779]= 16'h1df8;
assign q[8780]= 16'h18f8;
assign q[8781]= 16'h139b;
assign q[8782]= 16'hdf8;
assign q[8783]= 16'h825;
assign q[8784]= 16'h23d;
assign q[8785]= 16'hfc59;
assign q[8786]= 16'hf692;
assign q[8787]= 16'hf0ff;
assign q[8788]= 16'hebb9;
assign q[8789]= 16'he6d4;
assign q[8790]= 16'he263;
assign q[8791]= 16'hde76;
assign q[8792]= 16'hdb19;
assign q[8793]= 16'hd857;
assign q[8794]= 16'hd634;
assign q[8795]= 16'hd4b5;
assign q[8796]= 16'hd3d9;
assign q[8797]= 16'hd39d;
assign q[8798]= 16'hd3fc;
assign q[8799]= 16'hd4ee;
assign q[8800]= 16'hd668;
assign q[8801]= 16'hd85f;
assign q[8802]= 16'hdac5;
assign q[8803]= 16'hdd8d;
assign q[8804]= 16'he0a7;
assign q[8805]= 16'he402;
assign q[8806]= 16'he78f;
assign q[8807]= 16'heb3e;
assign q[8808]= 16'heeff;
assign q[8809]= 16'hf2c1;
assign q[8810]= 16'hf675;
assign q[8811]= 16'hfa0c;
assign q[8812]= 16'hfd79;
assign q[8813]= 16'hac;
assign q[8814]= 16'h39d;
assign q[8815]= 16'h63f;
assign q[8816]= 16'h889;
assign q[8817]= 16'ha72;
assign q[8818]= 16'hbf5;
assign q[8819]= 16'hd0e;
assign q[8820]= 16'hdb9;
assign q[8821]= 16'hdf7;
assign q[8822]= 16'hdca;
assign q[8823]= 16'hd35;
assign q[8824]= 16'hc41;
assign q[8825]= 16'haf5;
assign q[8826]= 16'h95c;
assign q[8827]= 16'h783;
assign q[8828]= 16'h579;
assign q[8829]= 16'h34e;
assign q[8830]= 16'h112;
assign q[8831]= 16'hfed9;
assign q[8832]= 16'hfcb3;
assign q[8833]= 16'hfab2;
assign q[8834]= 16'hf8e7;
assign q[8835]= 16'hf762;
assign q[8836]= 16'hf633;
assign q[8837]= 16'hf565;
assign q[8838]= 16'hf502;
assign q[8839]= 16'hf512;
assign q[8840]= 16'hf59a;
assign q[8841]= 16'hf69c;
assign q[8842]= 16'hf816;
assign q[8843]= 16'hfa06;
assign q[8844]= 16'hfc63;
assign q[8845]= 16'hff26;
assign q[8846]= 16'h241;
assign q[8847]= 16'h5a9;
assign q[8848]= 16'h94e;
assign q[8849]= 16'hd20;
assign q[8850]= 16'h110f;
assign q[8851]= 16'h150a;
assign q[8852]= 16'h18ff;
assign q[8853]= 16'h1ce0;
assign q[8854]= 16'h209d;
assign q[8855]= 16'h2427;
assign q[8856]= 16'h2773;
assign q[8857]= 16'h2a75;
assign q[8858]= 16'h2d25;
assign q[8859]= 16'h2f7a;
assign q[8860]= 16'h3171;
assign q[8861]= 16'h3305;
assign q[8862]= 16'h3434;
assign q[8863]= 16'h34fe;
assign q[8864]= 16'h3563;
assign q[8865]= 16'h3567;
assign q[8866]= 16'h350d;
assign q[8867]= 16'h3459;
assign q[8868]= 16'h3351;
assign q[8869]= 16'h31fd;
assign q[8870]= 16'h3062;
assign q[8871]= 16'h2e8a;
assign q[8872]= 16'h2c7d;
assign q[8873]= 16'h2a44;
assign q[8874]= 16'h27e9;
assign q[8875]= 16'h2577;
assign q[8876]= 16'h22f8;
assign q[8877]= 16'h2078;
assign q[8878]= 16'h1e02;
assign q[8879]= 16'h1ba0;
assign q[8880]= 16'h195e;
assign q[8881]= 16'h1747;
assign q[8882]= 16'h1563;
assign q[8883]= 16'h13bb;
assign q[8884]= 16'h1256;
assign q[8885]= 16'h113a;
assign q[8886]= 16'h106a;
assign q[8887]= 16'hfe6;
assign q[8888]= 16'hfae;
assign q[8889]= 16'hfbc;
assign q[8890]= 16'h100a;
assign q[8891]= 16'h108e;
assign q[8892]= 16'h113c;
assign q[8893]= 16'h1204;
assign q[8894]= 16'h12d8;
assign q[8895]= 16'h13a3;
assign q[8896]= 16'h1454;
assign q[8897]= 16'h14d7;
assign q[8898]= 16'h1519;
assign q[8899]= 16'h1507;
assign q[8900]= 16'h1493;
assign q[8901]= 16'h13af;
assign q[8902]= 16'h1250;
assign q[8903]= 16'h1070;
assign q[8904]= 16'he0e;
assign q[8905]= 16'hb2b;
assign q[8906]= 16'h7d1;
assign q[8907]= 16'h40a;
assign q[8908]= 16'hffe9;
assign q[8909]= 16'hfb81;
assign q[8910]= 16'hf6eb;
assign q[8911]= 16'hf245;
assign q[8912]= 16'hedab;
assign q[8913]= 16'he93d;
assign q[8914]= 16'he519;
assign q[8915]= 16'he15e;
assign q[8916]= 16'hde28;
assign q[8917]= 16'hdb8f;
assign q[8918]= 16'hd9a8;
assign q[8919]= 16'hd882;
assign q[8920]= 16'hd826;
assign q[8921]= 16'hd898;
assign q[8922]= 16'hd9d6;
assign q[8923]= 16'hdbd6;
assign q[8924]= 16'hde88;
assign q[8925]= 16'he1d6;
assign q[8926]= 16'he5a6;
assign q[8927]= 16'he9da;
assign q[8928]= 16'hee4f;
assign q[8929]= 16'hf2e2;
assign q[8930]= 16'hf76d;
assign q[8931]= 16'hfbcc;
assign q[8932]= 16'hffdf;
assign q[8933]= 16'h384;
assign q[8934]= 16'h6a3;
assign q[8935]= 16'h925;
assign q[8936]= 16'hafb;
assign q[8937]= 16'hc1d;
assign q[8938]= 16'hc87;
assign q[8939]= 16'hc40;
assign q[8940]= 16'hb53;
assign q[8941]= 16'h9d1;
assign q[8942]= 16'h7d3;
assign q[8943]= 16'h573;
assign q[8944]= 16'h2d3;
assign q[8945]= 16'h13;
assign q[8946]= 16'hfd58;
assign q[8947]= 16'hfac2;
assign q[8948]= 16'hf873;
assign q[8949]= 16'hf689;
assign q[8950]= 16'hf520;
assign q[8951]= 16'hf44b;
assign q[8952]= 16'hf41c;
assign q[8953]= 16'hf49b;
assign q[8954]= 16'hf5cd;
assign q[8955]= 16'hf7ad;
assign q[8956]= 16'hfa33;
assign q[8957]= 16'hfd4f;
assign q[8958]= 16'hec;
assign q[8959]= 16'h4f2;
assign q[8960]= 16'h944;
assign q[8961]= 16'hdc4;
assign q[8962]= 16'h1252;
assign q[8963]= 16'h16cd;
assign q[8964]= 16'h1b16;
assign q[8965]= 16'h1f12;
assign q[8966]= 16'h22a5;
assign q[8967]= 16'h25ba;
assign q[8968]= 16'h283f;
assign q[8969]= 16'h2a28;
assign q[8970]= 16'h2b6c;
assign q[8971]= 16'h2c0a;
assign q[8972]= 16'h2c05;
assign q[8973]= 16'h2b64;
assign q[8974]= 16'h2a32;
assign q[8975]= 16'h2881;
assign q[8976]= 16'h2661;
assign q[8977]= 16'h23e8;
assign q[8978]= 16'h212d;
assign q[8979]= 16'h1e46;
assign q[8980]= 16'h1b4a;
assign q[8981]= 16'h184f;
assign q[8982]= 16'h1569;
assign q[8983]= 16'h12aa;
assign q[8984]= 16'h1023;
assign q[8985]= 16'hde0;
assign q[8986]= 16'hbeb;
assign q[8987]= 16'ha4c;
assign q[8988]= 16'h907;
assign q[8989]= 16'h81c;
assign q[8990]= 16'h78d;
assign q[8991]= 16'h754;
assign q[8992]= 16'h76d;
assign q[8993]= 16'h7d3;
assign q[8994]= 16'h87e;
assign q[8995]= 16'h965;
assign q[8996]= 16'ha82;
assign q[8997]= 16'hbcb;
assign q[8998]= 16'hd3b;
assign q[8999]= 16'hec9;
assign q[9000]= 16'h106f;
assign q[9001]= 16'h1227;
assign q[9002]= 16'h13ec;
assign q[9003]= 16'h15ba;
assign q[9004]= 16'h178b;
assign q[9005]= 16'h195e;
assign q[9006]= 16'h1b2d;
assign q[9007]= 16'h1cf5;
assign q[9008]= 16'h1eb2;
assign q[9009]= 16'h2060;
assign q[9010]= 16'h21fb;
assign q[9011]= 16'h237e;
assign q[9012]= 16'h24e3;
assign q[9013]= 16'h2625;
assign q[9014]= 16'h273e;
assign q[9015]= 16'h2827;
assign q[9016]= 16'h28da;
assign q[9017]= 16'h2952;
assign q[9018]= 16'h2989;
assign q[9019]= 16'h297a;
assign q[9020]= 16'h2920;
assign q[9021]= 16'h287a;
assign q[9022]= 16'h2783;
assign q[9023]= 16'h263d;
assign q[9024]= 16'h24a7;
assign q[9025]= 16'h22c3;
assign q[9026]= 16'h2095;
assign q[9027]= 16'h1e20;
assign q[9028]= 16'h1b6b;
assign q[9029]= 16'h187d;
assign q[9030]= 16'h155b;
assign q[9031]= 16'h120f;
assign q[9032]= 16'hea0;
assign q[9033]= 16'hb15;
assign q[9034]= 16'h778;
assign q[9035]= 16'h3cf;
assign q[9036]= 16'h21;
assign q[9037]= 16'hfc76;
assign q[9038]= 16'hf8d0;
assign q[9039]= 16'hf536;
assign q[9040]= 16'hf1ac;
assign q[9041]= 16'hee34;
assign q[9042]= 16'head1;
assign q[9043]= 16'he785;
assign q[9044]= 16'he454;
assign q[9045]= 16'he13d;
assign q[9046]= 16'hde45;
assign q[9047]= 16'hdb6e;
assign q[9048]= 16'hd8bb;
assign q[9049]= 16'hd630;
assign q[9050]= 16'hd3d2;
assign q[9051]= 16'hd1a6;
assign q[9052]= 16'hcfb4;
assign q[9053]= 16'hce03;
assign q[9054]= 16'hcc9a;
assign q[9055]= 16'hcb82;
assign q[9056]= 16'hcac3;
assign q[9057]= 16'hca64;
assign q[9058]= 16'hca6d;
assign q[9059]= 16'hcae5;
assign q[9060]= 16'hcbcf;
assign q[9061]= 16'hcd2f;
assign q[9062]= 16'hcf05;
assign q[9063]= 16'hd150;
assign q[9064]= 16'hd40b;
assign q[9065]= 16'hd72e;
assign q[9066]= 16'hdab0;
assign q[9067]= 16'hde84;
assign q[9068]= 16'he299;
assign q[9069]= 16'he6dd;
assign q[9070]= 16'heb3e;
assign q[9071]= 16'hefa5;
assign q[9072]= 16'hf3fc;
assign q[9073]= 16'hf82d;
assign q[9074]= 16'hfc22;
assign q[9075]= 16'hffc4;
assign q[9076]= 16'h301;
assign q[9077]= 16'h5ca;
assign q[9078]= 16'h80f;
assign q[9079]= 16'h9c7;
assign q[9080]= 16'haec;
assign q[9081]= 16'hb7b;
assign q[9082]= 16'hb77;
assign q[9083]= 16'hae7;
assign q[9084]= 16'h9d7;
assign q[9085]= 16'h855;
assign q[9086]= 16'h674;
assign q[9087]= 16'h449;
assign q[9088]= 16'h1ec;
assign q[9089]= 16'hff77;
assign q[9090]= 16'hfd01;
assign q[9091]= 16'hfaa5;
assign q[9092]= 16'hf87b;
assign q[9093]= 16'hf698;
assign q[9094]= 16'hf510;
assign q[9095]= 16'hf3f1;
assign q[9096]= 16'hf349;
assign q[9097]= 16'hf31c;
assign q[9098]= 16'hf36d;
assign q[9099]= 16'hf43a;
assign q[9100]= 16'hf57c;
assign q[9101]= 16'hf725;
assign q[9102]= 16'hf927;
assign q[9103]= 16'hfb6d;
assign q[9104]= 16'hfde3;
assign q[9105]= 16'h6e;
assign q[9106]= 16'h2fa;
assign q[9107]= 16'h56b;
assign q[9108]= 16'h7ab;
assign q[9109]= 16'h9a3;
assign q[9110]= 16'hb41;
assign q[9111]= 16'hc76;
assign q[9112]= 16'hd34;
assign q[9113]= 16'hd77;
assign q[9114]= 16'hd39;
assign q[9115]= 16'hc7f;
assign q[9116]= 16'hb4f;
assign q[9117]= 16'h9b4;
assign q[9118]= 16'h7bd;
assign q[9119]= 16'h57c;
assign q[9120]= 16'h305;
assign q[9121]= 16'h6e;
assign q[9122]= 16'hfdcf;
assign q[9123]= 16'hfb3c;
assign q[9124]= 16'hf8cb;
assign q[9125]= 16'hf68e;
assign q[9126]= 16'hf497;
assign q[9127]= 16'hf2f0;
assign q[9128]= 16'hf1a4;
assign q[9129]= 16'hf0b5;
assign q[9130]= 16'hf023;
assign q[9131]= 16'hefea;
assign q[9132]= 16'hf001;
assign q[9133]= 16'hf05c;
assign q[9134]= 16'hf0e9;
assign q[9135]= 16'hf198;
assign q[9136]= 16'hf255;
assign q[9137]= 16'hf30a;
assign q[9138]= 16'hf3a4;
assign q[9139]= 16'hf410;
assign q[9140]= 16'hf43b;
assign q[9141]= 16'hf419;
assign q[9142]= 16'hf39e;
assign q[9143]= 16'hf2c3;
assign q[9144]= 16'hf186;
assign q[9145]= 16'hefe9;
assign q[9146]= 16'hedf3;
assign q[9147]= 16'hebaf;
assign q[9148]= 16'he92c;
assign q[9149]= 16'he67f;
assign q[9150]= 16'he3bc;
assign q[9151]= 16'he0fc;
assign q[9152]= 16'hde58;
assign q[9153]= 16'hdbea;
assign q[9154]= 16'hd9cc;
assign q[9155]= 16'hd815;
assign q[9156]= 16'hd6dc;
assign q[9157]= 16'hd633;
assign q[9158]= 16'hd629;
assign q[9159]= 16'hd6ca;
assign q[9160]= 16'hd81b;
assign q[9161]= 16'hda1f;
assign q[9162]= 16'hdcd3;
assign q[9163]= 16'he030;
assign q[9164]= 16'he42a;
assign q[9165]= 16'he8b1;
assign q[9166]= 16'hedb2;
assign q[9167]= 16'hf319;
assign q[9168]= 16'hf8cd;
assign q[9169]= 16'hfeb6;
assign q[9170]= 16'h4b8;
assign q[9171]= 16'habd;
assign q[9172]= 16'h10aa;
assign q[9173]= 16'h1668;
assign q[9174]= 16'h1be2;
assign q[9175]= 16'h2105;
assign q[9176]= 16'h25bf;
assign q[9177]= 16'h2a02;
assign q[9178]= 16'h2dc4;
assign q[9179]= 16'h30fc;
assign q[9180]= 16'h33a4;
assign q[9181]= 16'h35bb;
assign q[9182]= 16'h3741;
assign q[9183]= 16'h3837;
assign q[9184]= 16'h38a2;
assign q[9185]= 16'h3888;
assign q[9186]= 16'h37f1;
assign q[9187]= 16'h36e6;
assign q[9188]= 16'h3572;
assign q[9189]= 16'h33a0;
assign q[9190]= 16'h317c;
assign q[9191]= 16'h2f12;
assign q[9192]= 16'h2c72;
assign q[9193]= 16'h29a7;
assign q[9194]= 16'h26c2;
assign q[9195]= 16'h23d0;
assign q[9196]= 16'h20e0;
assign q[9197]= 16'h1e02;
assign q[9198]= 16'h1b43;
assign q[9199]= 16'h18b4;
assign q[9200]= 16'h1661;
assign q[9201]= 16'h1457;
assign q[9202]= 16'h12a3;
assign q[9203]= 16'h114f;
assign q[9204]= 16'h1063;
assign q[9205]= 16'hfe6;
assign q[9206]= 16'hfda;
assign q[9207]= 16'h1041;
assign q[9208]= 16'h1119;
assign q[9209]= 16'h125a;
assign q[9210]= 16'h13fd;
assign q[9211]= 16'h15f5;
assign q[9212]= 16'h1831;
assign q[9213]= 16'h1aa0;
assign q[9214]= 16'h1d2b;
assign q[9215]= 16'h1fbc;
assign q[9216]= 16'h2238;
assign q[9217]= 16'h2488;
assign q[9218]= 16'h268f;
assign q[9219]= 16'h2837;
assign q[9220]= 16'h2966;
assign q[9221]= 16'h2a09;
assign q[9222]= 16'h2a0d;
assign q[9223]= 16'h2964;
assign q[9224]= 16'h2804;
assign q[9225]= 16'h25ea;
assign q[9226]= 16'h2316;
assign q[9227]= 16'h1f8d;
assign q[9228]= 16'h1b5b;
assign q[9229]= 16'h1691;
assign q[9230]= 16'h1142;
assign q[9231]= 16'hb89;
assign q[9232]= 16'h581;
assign q[9233]= 16'hff4a;
assign q[9234]= 16'hf902;
assign q[9235]= 16'hf2ca;
assign q[9236]= 16'hecc1;
assign q[9237]= 16'he705;
assign q[9238]= 16'he1b2;
assign q[9239]= 16'hdcde;
assign q[9240]= 16'hd89d;
assign q[9241]= 16'hd4fc;
assign q[9242]= 16'hd204;
assign q[9243]= 16'hcfb8;
assign q[9244]= 16'hce14;
assign q[9245]= 16'hcd12;
assign q[9246]= 16'hcca3;
assign q[9247]= 16'hccb6;
assign q[9248]= 16'hcd36;
assign q[9249]= 16'hce0c;
assign q[9250]= 16'hcf1e;
assign q[9251]= 16'hd053;
assign q[9252]= 16'hd191;
assign q[9253]= 16'hd2c1;
assign q[9254]= 16'hd3ce;
assign q[9255]= 16'hd4a6;
assign q[9256]= 16'hd53d;
assign q[9257]= 16'hd58b;
assign q[9258]= 16'hd58b;
assign q[9259]= 16'hd53f;
assign q[9260]= 16'hd4b0;
assign q[9261]= 16'hd3e8;
assign q[9262]= 16'hd2f7;
assign q[9263]= 16'hd1f2;
assign q[9264]= 16'hd0ed;
assign q[9265]= 16'hd002;
assign q[9266]= 16'hcf47;
assign q[9267]= 16'hced5;
assign q[9268]= 16'hcec2;
assign q[9269]= 16'hcf21;
assign q[9270]= 16'hd001;
assign q[9271]= 16'hd16c;
assign q[9272]= 16'hd36a;
assign q[9273]= 16'hd5f9;
assign q[9274]= 16'hd914;
assign q[9275]= 16'hdcb0;
assign q[9276]= 16'he0bc;
assign q[9277]= 16'he520;
assign q[9278]= 16'he9c4;
assign q[9279]= 16'hee88;
assign q[9280]= 16'hf34d;
assign q[9281]= 16'hf7f1;
assign q[9282]= 16'hfc52;
assign q[9283]= 16'h4e;
assign q[9284]= 16'h3c9;
assign q[9285]= 16'h6a8;
assign q[9286]= 16'h8d3;
assign q[9287]= 16'ha3a;
assign q[9288]= 16'had2;
assign q[9289]= 16'ha96;
assign q[9290]= 16'h989;
assign q[9291]= 16'h7b3;
assign q[9292]= 16'h522;
assign q[9293]= 16'h1ed;
assign q[9294]= 16'hfe2e;
assign q[9295]= 16'hfa02;
assign q[9296]= 16'hf58a;
assign q[9297]= 16'hf0e9;
assign q[9298]= 16'hec45;
assign q[9299]= 16'he7c1;
assign q[9300]= 16'he37e;
assign q[9301]= 16'hdf9b;
assign q[9302]= 16'hdc34;
assign q[9303]= 16'hd95f;
assign q[9304]= 16'hd72c;
assign q[9305]= 16'hd5a6;
assign q[9306]= 16'hd4d2;
assign q[9307]= 16'hd4ae;
assign q[9308]= 16'hd533;
assign q[9309]= 16'hd654;
assign q[9310]= 16'hd7ff;
assign q[9311]= 16'hda1d;
assign q[9312]= 16'hdc97;
assign q[9313]= 16'hdf50;
assign q[9314]= 16'he22d;
assign q[9315]= 16'he512;
assign q[9316]= 16'he7e4;
assign q[9317]= 16'hea8c;
assign q[9318]= 16'hecf3;
assign q[9319]= 16'hef0a;
assign q[9320]= 16'hf0c3;
assign q[9321]= 16'hf216;
assign q[9322]= 16'hf302;
assign q[9323]= 16'hf389;
assign q[9324]= 16'hf3b1;
assign q[9325]= 16'hf386;
assign q[9326]= 16'hf318;
assign q[9327]= 16'hf278;
assign q[9328]= 16'hf1bb;
assign q[9329]= 16'hf0f5;
assign q[9330]= 16'hf03c;
assign q[9331]= 16'hefa6;
assign q[9332]= 16'hef43;
assign q[9333]= 16'hef25;
assign q[9334]= 16'hef58;
assign q[9335]= 16'hefe5;
assign q[9336]= 16'hf0d1;
assign q[9337]= 16'hf21c;
assign q[9338]= 16'hf3c1;
assign q[9339]= 16'hf5b9;
assign q[9340]= 16'hf7f5;
assign q[9341]= 16'hfa66;
assign q[9342]= 16'hfcf9;
assign q[9343]= 16'hff97;
assign q[9344]= 16'h22a;
assign q[9345]= 16'h49d;
assign q[9346]= 16'h6d7;
assign q[9347]= 16'h8c3;
assign q[9348]= 16'ha4e;
assign q[9349]= 16'hb67;
assign q[9350]= 16'hc02;
assign q[9351]= 16'hc13;
assign q[9352]= 16'hb96;
assign q[9353]= 16'ha8a;
assign q[9354]= 16'h8f0;
assign q[9355]= 16'h6d1;
assign q[9356]= 16'h436;
assign q[9357]= 16'h12d;
assign q[9358]= 16'hfdc7;
assign q[9359]= 16'hfa15;
assign q[9360]= 16'hf62b;
assign q[9361]= 16'hf21e;
assign q[9362]= 16'hee02;
assign q[9363]= 16'he9ec;
assign q[9364]= 16'he5ed;
assign q[9365]= 16'he217;
assign q[9366]= 16'hde7a;
assign q[9367]= 16'hdb22;
assign q[9368]= 16'hd81a;
assign q[9369]= 16'hd569;
assign q[9370]= 16'hd314;
assign q[9371]= 16'hd11f;
assign q[9372]= 16'hcf89;
assign q[9373]= 16'hce51;
assign q[9374]= 16'hcd73;
assign q[9375]= 16'hcceb;
assign q[9376]= 16'hccb2;
assign q[9377]= 16'hccc1;
assign q[9378]= 16'hcd10;
assign q[9379]= 16'hcd98;
assign q[9380]= 16'hce50;
assign q[9381]= 16'hcf2f;
assign q[9382]= 16'hd02d;
assign q[9383]= 16'hd143;
assign q[9384]= 16'hd266;
assign q[9385]= 16'hd391;
assign q[9386]= 16'hd4b9;
assign q[9387]= 16'hd5d8;
assign q[9388]= 16'hd6e5;
assign q[9389]= 16'hd7d9;
assign q[9390]= 16'hd8ac;
assign q[9391]= 16'hd957;
assign q[9392]= 16'hd9d3;
assign q[9393]= 16'hda19;
assign q[9394]= 16'hda25;
assign q[9395]= 16'hd9f3;
assign q[9396]= 16'hd97f;
assign q[9397]= 16'hd8ca;
assign q[9398]= 16'hd7d4;
assign q[9399]= 16'hd6a3;
assign q[9400]= 16'hd53b;
assign q[9401]= 16'hd3a7;
assign q[9402]= 16'hd1f2;
assign q[9403]= 16'hd02a;
assign q[9404]= 16'hce61;
assign q[9405]= 16'hccab;
assign q[9406]= 16'hcb1b;
assign q[9407]= 16'hc9c8;
assign q[9408]= 16'hc8c7;
assign q[9409]= 16'hc831;
assign q[9410]= 16'hc818;
assign q[9411]= 16'hc890;
assign q[9412]= 16'hc9aa;
assign q[9413]= 16'hcb71;
assign q[9414]= 16'hcdee;
assign q[9415]= 16'hd123;
assign q[9416]= 16'hd50f;
assign q[9417]= 16'hd9a8;
assign q[9418]= 16'hdee0;
assign q[9419]= 16'he4a4;
assign q[9420]= 16'head9;
assign q[9421]= 16'hf161;
assign q[9422]= 16'hf819;
assign q[9423]= 16'hfedb;
assign q[9424]= 16'h57e;
assign q[9425]= 16'hbd9;
assign q[9426]= 16'h11c5;
assign q[9427]= 16'h1718;
assign q[9428]= 16'h1baf;
assign q[9429]= 16'h1f6b;
assign q[9430]= 16'h2230;
assign q[9431]= 16'h23ea;
assign q[9432]= 16'h248e;
assign q[9433]= 16'h2416;
assign q[9434]= 16'h2285;
assign q[9435]= 16'h1fe7;
assign q[9436]= 16'h1c4f;
assign q[9437]= 16'h17d8;
assign q[9438]= 16'h12a4;
assign q[9439]= 16'hcd8;
assign q[9440]= 16'h6a0;
assign q[9441]= 16'h2a;
assign q[9442]= 16'hf9a7;
assign q[9443]= 16'hf344;
assign q[9444]= 16'hed30;
assign q[9445]= 16'he797;
assign q[9446]= 16'he29f;
assign q[9447]= 16'hde69;
assign q[9448]= 16'hdb11;
assign q[9449]= 16'hd8ab;
assign q[9450]= 16'hd743;
assign q[9451]= 16'hd6de;
assign q[9452]= 16'hd779;
assign q[9453]= 16'hd90a;
assign q[9454]= 16'hdb80;
assign q[9455]= 16'hdec5;
assign q[9456]= 16'he2be;
assign q[9457]= 16'he74b;
assign q[9458]= 16'hec4c;
assign q[9459]= 16'hf19e;
assign q[9460]= 16'hf71e;
assign q[9461]= 16'hfcab;
assign q[9462]= 16'h224;
assign q[9463]= 16'h770;
assign q[9464]= 16'hc76;
assign q[9465]= 16'h1122;
assign q[9466]= 16'h1564;
assign q[9467]= 16'h1932;
assign q[9468]= 16'h1c88;
assign q[9469]= 16'h1f64;
assign q[9470]= 16'h21ca;
assign q[9471]= 16'h23c0;
assign q[9472]= 16'h254f;
assign q[9473]= 16'h2685;
assign q[9474]= 16'h276d;
assign q[9475]= 16'h2816;
assign q[9476]= 16'h288e;
assign q[9477]= 16'h28e1;
assign q[9478]= 16'h291b;
assign q[9479]= 16'h2948;
assign q[9480]= 16'h296f;
assign q[9481]= 16'h2997;
assign q[9482]= 16'h29c3;
assign q[9483]= 16'h29f8;
assign q[9484]= 16'h2a34;
assign q[9485]= 16'h2a78;
assign q[9486]= 16'h2ac1;
assign q[9487]= 16'h2b0d;
assign q[9488]= 16'h2b58;
assign q[9489]= 16'h2ba0;
assign q[9490]= 16'h2be2;
assign q[9491]= 16'h2c1c;
assign q[9492]= 16'h2c4c;
assign q[9493]= 16'h2c71;
assign q[9494]= 16'h2c8d;
assign q[9495]= 16'h2ca0;
assign q[9496]= 16'h2cad;
assign q[9497]= 16'h2cb5;
assign q[9498]= 16'h2cbc;
assign q[9499]= 16'h2cc4;
assign q[9500]= 16'h2ccf;
assign q[9501]= 16'h2cdf;
assign q[9502]= 16'h2cf5;
assign q[9503]= 16'h2d11;
assign q[9504]= 16'h2d32;
assign q[9505]= 16'h2d57;
assign q[9506]= 16'h2d7b;
assign q[9507]= 16'h2d9c;
assign q[9508]= 16'h2db5;
assign q[9509]= 16'h2dc2;
assign q[9510]= 16'h2dbe;
assign q[9511]= 16'h2da5;
assign q[9512]= 16'h2d74;
assign q[9513]= 16'h2d29;
assign q[9514]= 16'h2cc4;
assign q[9515]= 16'h2c46;
assign q[9516]= 16'h2bb2;
assign q[9517]= 16'h2b0e;
assign q[9518]= 16'h2a61;
assign q[9519]= 16'h29b3;
assign q[9520]= 16'h290e;
assign q[9521]= 16'h287e;
assign q[9522]= 16'h280d;
assign q[9523]= 16'h27c7;
assign q[9524]= 16'h27b5;
assign q[9525]= 16'h27df;
assign q[9526]= 16'h284c;
assign q[9527]= 16'h28ff;
assign q[9528]= 16'h29f6;
assign q[9529]= 16'h2b2f;
assign q[9530]= 16'h2ca0;
assign q[9531]= 16'h2e3e;
assign q[9532]= 16'h2ff8;
assign q[9533]= 16'h31ba;
assign q[9534]= 16'h336e;
assign q[9535]= 16'h34f9;
assign q[9536]= 16'h3642;
assign q[9537]= 16'h372d;
assign q[9538]= 16'h379f;
assign q[9539]= 16'h3781;
assign q[9540]= 16'h36bb;
assign q[9541]= 16'h353d;
assign q[9542]= 16'h32fa;
assign q[9543]= 16'h2feb;
assign q[9544]= 16'h2c11;
assign q[9545]= 16'h2773;
assign q[9546]= 16'h221e;
assign q[9547]= 16'h1c2a;
assign q[9548]= 16'h15b2;
assign q[9549]= 16'hed8;
assign q[9550]= 16'h7c4;
assign q[9551]= 16'ha3;
assign q[9552]= 16'hf9a3;
assign q[9553]= 16'hf2f1;
assign q[9554]= 16'hecbe;
assign q[9555]= 16'he737;
assign q[9556]= 16'he283;
assign q[9557]= 16'hdec7;
assign q[9558]= 16'hdc1f;
assign q[9559]= 16'hdaa1;
assign q[9560]= 16'hda57;
assign q[9561]= 16'hdb45;
assign q[9562]= 16'hdd62;
assign q[9563]= 16'he09f;
assign q[9564]= 16'he4e0;
assign q[9565]= 16'hea03;
assign q[9566]= 16'hefdd;
assign q[9567]= 16'hf63e;
assign q[9568]= 16'hfcf1;
assign q[9569]= 16'h3bd;
assign q[9570]= 16'ha6c;
assign q[9571]= 16'h10c3;
assign q[9572]= 16'h168f;
assign q[9573]= 16'h1b9f;
assign q[9574]= 16'h1fc9;
assign q[9575]= 16'h22ea;
assign q[9576]= 16'h24e7;
assign q[9577]= 16'h25b1;
assign q[9578]= 16'h2541;
assign q[9579]= 16'h239a;
assign q[9580]= 16'h20c9;
assign q[9581]= 16'h1ce4;
assign q[9582]= 16'h1809;
assign q[9583]= 16'h125e;
assign q[9584]= 16'hc0d;
assign q[9585]= 16'h545;
assign q[9586]= 16'hfe37;
assign q[9587]= 16'hf713;
assign q[9588]= 16'hf009;
assign q[9589]= 16'he946;
assign q[9590]= 16'he2f2;
assign q[9591]= 16'hdd30;
assign q[9592]= 16'hd81d;
assign q[9593]= 16'hd3cb;
assign q[9594]= 16'hd049;
assign q[9595]= 16'hcd9a;
assign q[9596]= 16'hcbbb;
assign q[9597]= 16'hcaa2;
assign q[9598]= 16'hca3c;
assign q[9599]= 16'hca75;
assign q[9600]= 16'hcb30;
assign q[9601]= 16'hcc50;
assign q[9602]= 16'hcdb5;
assign q[9603]= 16'hcf3f;
assign q[9604]= 16'hd0d0;
assign q[9605]= 16'hd24d;
assign q[9606]= 16'hd39c;
assign q[9607]= 16'hd4a9;
assign q[9608]= 16'hd568;
assign q[9609]= 16'hd5cf;
assign q[9610]= 16'hd5dc;
assign q[9611]= 16'hd593;
assign q[9612]= 16'hd4fd;
assign q[9613]= 16'hd429;
assign q[9614]= 16'hd32a;
assign q[9615]= 16'hd217;
assign q[9616]= 16'hd109;
assign q[9617]= 16'hd01c;
assign q[9618]= 16'hcf69;
assign q[9619]= 16'hcf0c;
assign q[9620]= 16'hcf1c;
assign q[9621]= 16'hcfae;
assign q[9622]= 16'hd0d3;
assign q[9623]= 16'hd297;
assign q[9624]= 16'hd501;
assign q[9625]= 16'hd813;
assign q[9626]= 16'hdbc9;
assign q[9627]= 16'he01a;
assign q[9628]= 16'he4f7;
assign q[9629]= 16'hea4d;
assign q[9630]= 16'hf005;
assign q[9631]= 16'hf605;
assign q[9632]= 16'hfc2f;
assign q[9633]= 16'h266;
assign q[9634]= 16'h88d;
assign q[9635]= 16'he86;
assign q[9636]= 16'h1433;
assign q[9637]= 16'h197b;
assign q[9638]= 16'h1e47;
assign q[9639]= 16'h2283;
assign q[9640]= 16'h261f;
assign q[9641]= 16'h290f;
assign q[9642]= 16'h2b4d;
assign q[9643]= 16'h2cd4;
assign q[9644]= 16'h2da6;
assign q[9645]= 16'h2dc5;
assign q[9646]= 16'h2d3b;
assign q[9647]= 16'h2c12;
assign q[9648]= 16'h2a55;
assign q[9649]= 16'h2813;
assign q[9650]= 16'h255c;
assign q[9651]= 16'h2240;
assign q[9652]= 16'h1ecf;
assign q[9653]= 16'h1b17;
assign q[9654]= 16'h172a;
assign q[9655]= 16'h1315;
assign q[9656]= 16'hee4;
assign q[9657]= 16'haa4;
assign q[9658]= 16'h660;
assign q[9659]= 16'h221;
assign q[9660]= 16'hfdf0;
assign q[9661]= 16'hf9d2;
assign q[9662]= 16'hf5cf;
assign q[9663]= 16'hf1ed;
assign q[9664]= 16'hee31;
assign q[9665]= 16'hea9f;
assign q[9666]= 16'he73d;
assign q[9667]= 16'he40e;
assign q[9668]= 16'he117;
assign q[9669]= 16'hde5b;
assign q[9670]= 16'hdbde;
assign q[9671]= 16'hd9a3;
assign q[9672]= 16'hd7ac;
assign q[9673]= 16'hd5fb;
assign q[9674]= 16'hd490;
assign q[9675]= 16'hd36b;
assign q[9676]= 16'hd28a;
assign q[9677]= 16'hd1eb;
assign q[9678]= 16'hd188;
assign q[9679]= 16'hd15d;
assign q[9680]= 16'hd161;
assign q[9681]= 16'hd18e;
assign q[9682]= 16'hd1da;
assign q[9683]= 16'hd23b;
assign q[9684]= 16'hd2a9;
assign q[9685]= 16'hd318;
assign q[9686]= 16'hd380;
assign q[9687]= 16'hd3d8;
assign q[9688]= 16'hd41a;
assign q[9689]= 16'hd440;
assign q[9690]= 16'hd447;
assign q[9691]= 16'hd42e;
assign q[9692]= 16'hd3f6;
assign q[9693]= 16'hd3a2;
assign q[9694]= 16'hd338;
assign q[9695]= 16'hd2c0;
assign q[9696]= 16'hd243;
assign q[9697]= 16'hd1cc;
assign q[9698]= 16'hd167;
assign q[9699]= 16'hd121;
assign q[9700]= 16'hd105;
assign q[9701]= 16'hd11e;
assign q[9702]= 16'hd176;
assign q[9703]= 16'hd215;
assign q[9704]= 16'hd300;
assign q[9705]= 16'hd43a;
assign q[9706]= 16'hd5c1;
assign q[9707]= 16'hd792;
assign q[9708]= 16'hd9a5;
assign q[9709]= 16'hdbf0;
assign q[9710]= 16'hde66;
assign q[9711]= 16'he0f7;
assign q[9712]= 16'he391;
assign q[9713]= 16'he622;
assign q[9714]= 16'he898;
assign q[9715]= 16'headf;
assign q[9716]= 16'hece7;
assign q[9717]= 16'heea2;
assign q[9718]= 16'hf003;
assign q[9719]= 16'hf101;
assign q[9720]= 16'hf19a;
assign q[9721]= 16'hf1cd;
assign q[9722]= 16'hf19f;
assign q[9723]= 16'hf11b;
assign q[9724]= 16'hf04e;
assign q[9725]= 16'hef4b;
assign q[9726]= 16'hee27;
assign q[9727]= 16'hecfc;
assign q[9728]= 16'hebe3;
assign q[9729]= 16'heaf7;
assign q[9730]= 16'hea52;
assign q[9731]= 16'hea0e;
assign q[9732]= 16'hea41;
assign q[9733]= 16'heafe;
assign q[9734]= 16'hec50;
assign q[9735]= 16'hee42;
assign q[9736]= 16'hf0d5;
assign q[9737]= 16'hf405;
assign q[9738]= 16'hf7c6;
assign q[9739]= 16'hfc08;
assign q[9740]= 16'hb1;
assign q[9741]= 16'h5a7;
assign q[9742]= 16'hac7;
assign q[9743]= 16'hfec;
assign q[9744]= 16'h14ef;
assign q[9745]= 16'h19a8;
assign q[9746]= 16'h1df0;
assign q[9747]= 16'h21a1;
assign q[9748]= 16'h249a;
assign q[9749]= 16'h26bd;
assign q[9750]= 16'h27f3;
assign q[9751]= 16'h282d;
assign q[9752]= 16'h2761;
assign q[9753]= 16'h2590;
assign q[9754]= 16'h22c0;
assign q[9755]= 16'h1f03;
assign q[9756]= 16'h1a6e;
assign q[9757]= 16'h1523;
assign q[9758]= 16'hf43;
assign q[9759]= 16'h8fb;
assign q[9760]= 16'h275;
assign q[9761]= 16'hfbe3;
assign q[9762]= 16'hf572;
assign q[9763]= 16'hef50;
assign q[9764]= 16'he9a9;
assign q[9765]= 16'he4a4;
assign q[9766]= 16'he063;
assign q[9767]= 16'hdd02;
assign q[9768]= 16'hda94;
assign q[9769]= 16'hd925;
assign q[9770]= 16'hd8b8;
assign q[9771]= 16'hd94a;
assign q[9772]= 16'hdace;
assign q[9773]= 16'hdd30;
assign q[9774]= 16'he056;
assign q[9775]= 16'he420;
assign q[9776]= 16'he869;
assign q[9777]= 16'hed0b;
assign q[9778]= 16'hf1de;
assign q[9779]= 16'hf6b7;
assign q[9780]= 16'hfb71;
assign q[9781]= 16'hffe6;
assign q[9782]= 16'h3f3;
assign q[9783]= 16'h77e;
assign q[9784]= 16'ha6e;
assign q[9785]= 16'hcb4;
assign q[9786]= 16'he44;
assign q[9787]= 16'hf1a;
assign q[9788]= 16'hf38;
assign q[9789]= 16'hea7;
assign q[9790]= 16'hd74;
assign q[9791]= 16'hbb1;
assign q[9792]= 16'h974;
assign q[9793]= 16'h6d6;
assign q[9794]= 16'h3f2;
assign q[9795]= 16'he3;
assign q[9796]= 16'hfdc4;
assign q[9797]= 16'hfaad;
assign q[9798]= 16'hf7b7;
assign q[9799]= 16'hf4f7;
assign q[9800]= 16'hf27d;
assign q[9801]= 16'hf058;
assign q[9802]= 16'hee91;
assign q[9803]= 16'hed2c;
assign q[9804]= 16'hec2c;
assign q[9805]= 16'heb8d;
assign q[9806]= 16'heb4a;
assign q[9807]= 16'heb5a;
assign q[9808]= 16'hebb1;
assign q[9809]= 16'hec42;
assign q[9810]= 16'hecff;
assign q[9811]= 16'hedda;
assign q[9812]= 16'heec3;
assign q[9813]= 16'hefaf;
assign q[9814]= 16'hf08f;
assign q[9815]= 16'hf15b;
assign q[9816]= 16'hf209;
assign q[9817]= 16'hf293;
assign q[9818]= 16'hf2f6;
assign q[9819]= 16'hf330;
assign q[9820]= 16'hf343;
assign q[9821]= 16'hf331;
assign q[9822]= 16'hf300;
assign q[9823]= 16'hf2b7;
assign q[9824]= 16'hf25d;
assign q[9825]= 16'hf1fc;
assign q[9826]= 16'hf19c;
assign q[9827]= 16'hf147;
assign q[9828]= 16'hf107;
assign q[9829]= 16'hf0e3;
assign q[9830]= 16'hf0e4;
assign q[9831]= 16'hf110;
assign q[9832]= 16'hf16d;
assign q[9833]= 16'hf1fe;
assign q[9834]= 16'hf2c6;
assign q[9835]= 16'hf3c5;
assign q[9836]= 16'hf4fb;
assign q[9837]= 16'hf667;
assign q[9838]= 16'hf806;
assign q[9839]= 16'hf9d2;
assign q[9840]= 16'hfbc9;
assign q[9841]= 16'hfde3;
assign q[9842]= 16'h1a;
assign q[9843]= 16'h26a;
assign q[9844]= 16'h4cc;
assign q[9845]= 16'h739;
assign q[9846]= 16'h9ab;
assign q[9847]= 16'hc1c;
assign q[9848]= 16'he88;
assign q[9849]= 16'h10ea;
assign q[9850]= 16'h133d;
assign q[9851]= 16'h157d;
assign q[9852]= 16'h17a9;
assign q[9853]= 16'h19bc;
assign q[9854]= 16'h1bb5;
assign q[9855]= 16'h1d92;
assign q[9856]= 16'h1f51;
assign q[9857]= 16'h20f1;
assign q[9858]= 16'h2270;
assign q[9859]= 16'h23cd;
assign q[9860]= 16'h2506;
assign q[9861]= 16'h261a;
assign q[9862]= 16'h2705;
assign q[9863]= 16'h27c6;
assign q[9864]= 16'h285b;
assign q[9865]= 16'h28bf;
assign q[9866]= 16'h28ef;
assign q[9867]= 16'h28e9;
assign q[9868]= 16'h28a8;
assign q[9869]= 16'h2829;
assign q[9870]= 16'h2768;
assign q[9871]= 16'h2663;
assign q[9872]= 16'h2518;
assign q[9873]= 16'h2384;
assign q[9874]= 16'h21a7;
assign q[9875]= 16'h1f83;
assign q[9876]= 16'h1d18;
assign q[9877]= 16'h1a6c;
assign q[9878]= 16'h1784;
assign q[9879]= 16'h1467;
assign q[9880]= 16'h111e;
assign q[9881]= 16'hdb5;
assign q[9882]= 16'ha39;
assign q[9883]= 16'h6b8;
assign q[9884]= 16'h342;
assign q[9885]= 16'hffe9;
assign q[9886]= 16'hfcbd;
assign q[9887]= 16'hf9d1;
assign q[9888]= 16'hf736;
assign q[9889]= 16'hf4fe;
assign q[9890]= 16'hf338;
assign q[9891]= 16'hf1f2;
assign q[9892]= 16'hf137;
assign q[9893]= 16'hf10f;
assign q[9894]= 16'hf181;
assign q[9895]= 16'hf28e;
assign q[9896]= 16'hf433;
assign q[9897]= 16'hf66b;
assign q[9898]= 16'hf92a;
assign q[9899]= 16'hfc63;
assign q[9900]= 16'h2;
assign q[9901]= 16'h3f4;
assign q[9902]= 16'h81f;
assign q[9903]= 16'hc69;
assign q[9904]= 16'h10b6;
assign q[9905]= 16'h14e8;
assign q[9906]= 16'h18e2;
assign q[9907]= 16'h1c8a;
assign q[9908]= 16'h1fc3;
assign q[9909]= 16'h2278;
assign q[9910]= 16'h2493;
assign q[9911]= 16'h2605;
assign q[9912]= 16'h26c2;
assign q[9913]= 16'h26c5;
assign q[9914]= 16'h260b;
assign q[9915]= 16'h249a;
assign q[9916]= 16'h227b;
assign q[9917]= 16'h1fbd;
assign q[9918]= 16'h1c75;
assign q[9919]= 16'h18b8;
assign q[9920]= 16'h14a3;
assign q[9921]= 16'h1053;
assign q[9922]= 16'hbe7;
assign q[9923]= 16'h77d;
assign q[9924]= 16'h337;
assign q[9925]= 16'hff30;
assign q[9926]= 16'hfb85;
assign q[9927]= 16'hf84c;
assign q[9928]= 16'hf59b;
assign q[9929]= 16'hf382;
assign q[9930]= 16'hf20a;
assign q[9931]= 16'hf13b;
assign q[9932]= 16'hf114;
assign q[9933]= 16'hf191;
assign q[9934]= 16'hf2a9;
assign q[9935]= 16'hf44f;
assign q[9936]= 16'hf672;
assign q[9937]= 16'hf8fd;
assign q[9938]= 16'hfbdc;
assign q[9939]= 16'hfef8;
assign q[9940]= 16'h239;
assign q[9941]= 16'h589;
assign q[9942]= 16'h8d5;
assign q[9943]= 16'hc08;
assign q[9944]= 16'hf14;
assign q[9945]= 16'h11eb;
assign q[9946]= 16'h1485;
assign q[9947]= 16'h16dd;
assign q[9948]= 16'h18f2;
assign q[9949]= 16'h1ac6;
assign q[9950]= 16'h1c5f;
assign q[9951]= 16'h1dc4;
assign q[9952]= 16'h1f00;
assign q[9953]= 16'h201f;
assign q[9954]= 16'h212d;
assign q[9955]= 16'h2237;
assign q[9956]= 16'h2346;
assign q[9957]= 16'h2466;
assign q[9958]= 16'h259e;
assign q[9959]= 16'h26f1;
assign q[9960]= 16'h2863;
assign q[9961]= 16'h29f0;
assign q[9962]= 16'h2b93;
assign q[9963]= 16'h2d43;
assign q[9964]= 16'h2ef4;
assign q[9965]= 16'h3096;
assign q[9966]= 16'h321a;
assign q[9967]= 16'h336b;
assign q[9968]= 16'h3476;
assign q[9969]= 16'h3527;
assign q[9970]= 16'h356c;
assign q[9971]= 16'h3533;
assign q[9972]= 16'h346d;
assign q[9973]= 16'h330f;
assign q[9974]= 16'h3110;
assign q[9975]= 16'h2e6d;
assign q[9976]= 16'h2b26;
assign q[9977]= 16'h2741;
assign q[9978]= 16'h22c9;
assign q[9979]= 16'h1dcc;
assign q[9980]= 16'h185d;
assign q[9981]= 16'h1292;
assign q[9982]= 16'hc86;
assign q[9983]= 16'h653;
assign q[9984]= 16'h18;
assign q[9985]= 16'hf9f3;
assign q[9986]= 16'hf400;
assign q[9987]= 16'hee5b;
assign q[9988]= 16'he920;
assign q[9989]= 16'he465;
assign q[9990]= 16'he03d;
assign q[9991]= 16'hdcb9;
assign q[9992]= 16'hd9e3;
assign q[9993]= 16'hd7c1;
assign q[9994]= 16'hd655;
assign q[9995]= 16'hd59c;
assign q[9996]= 16'hd58e;
assign q[9997]= 16'hd61e;
assign q[9998]= 16'hd73e;
assign q[9999]= 16'hd8db;
assign q[10000]= 16'hdadf;
assign q[10001]= 16'hdd36;
assign q[10002]= 16'hdfc7;
assign q[10003]= 16'he27b;
assign q[10004]= 16'he53c;
assign q[10005]= 16'he7f4;
assign q[10006]= 16'hea91;
assign q[10007]= 16'hed02;
assign q[10008]= 16'hef39;
assign q[10009]= 16'hf12a;
assign q[10010]= 16'hf2cf;
assign q[10011]= 16'hf422;
assign q[10012]= 16'hf523;
assign q[10013]= 16'hf5d3;
assign q[10014]= 16'hf636;
assign q[10015]= 16'hf652;
assign q[10016]= 16'hf630;
assign q[10017]= 16'hf5d9;
assign q[10018]= 16'hf558;
assign q[10019]= 16'hf4b6;
assign q[10020]= 16'hf400;
assign q[10021]= 16'hf33e;
assign q[10022]= 16'hf27b;
assign q[10023]= 16'hf1bf;
assign q[10024]= 16'hf111;
assign q[10025]= 16'hf077;
assign q[10026]= 16'heff4;
assign q[10027]= 16'hef8b;
assign q[10028]= 16'hef3f;
assign q[10029]= 16'hef0e;
assign q[10030]= 16'heef8;
assign q[10031]= 16'heefa;
assign q[10032]= 16'hef12;
assign q[10033]= 16'hef3d;
assign q[10034]= 16'hef77;
assign q[10035]= 16'hefbc;
assign q[10036]= 16'hf009;
assign q[10037]= 16'hf05c;
assign q[10038]= 16'hf0af;
assign q[10039]= 16'hf102;
assign q[10040]= 16'hf152;
assign q[10041]= 16'hf19d;
assign q[10042]= 16'hf1e2;
assign q[10043]= 16'hf21f;
assign q[10044]= 16'hf254;
assign q[10045]= 16'hf280;
assign q[10046]= 16'hf2a2;
assign q[10047]= 16'hf2ba;
assign q[10048]= 16'hf2c8;
assign q[10049]= 16'hf2ca;
assign q[10050]= 16'hf2c0;
assign q[10051]= 16'hf2ab;
assign q[10052]= 16'hf288;
assign q[10053]= 16'hf25a;
assign q[10054]= 16'hf21e;
assign q[10055]= 16'hf1d7;
assign q[10056]= 16'hf184;
assign q[10057]= 16'hf127;
assign q[10058]= 16'hf0c3;
assign q[10059]= 16'hf059;
assign q[10060]= 16'hefee;
assign q[10061]= 16'hef86;
assign q[10062]= 16'hef25;
assign q[10063]= 16'heed1;
assign q[10064]= 16'hee8f;
assign q[10065]= 16'hee65;
assign q[10066]= 16'hee5a;
assign q[10067]= 16'hee72;
assign q[10068]= 16'heeb4;
assign q[10069]= 16'hef23;
assign q[10070]= 16'hefc4;
assign q[10071]= 16'hf098;
assign q[10072]= 16'hf1a0;
assign q[10073]= 16'hf2dd;
assign q[10074]= 16'hf44c;
assign q[10075]= 16'hf5ea;
assign q[10076]= 16'hf7b1;
assign q[10077]= 16'hf99b;
assign q[10078]= 16'hfba0;
assign q[10079]= 16'hfdb7;
assign q[10080]= 16'hffd6;
assign q[10081]= 16'h1f2;
assign q[10082]= 16'h402;
assign q[10083]= 16'h5fd;
assign q[10084]= 16'h7d8;
assign q[10085]= 16'h98b;
assign q[10086]= 16'hb0f;
assign q[10087]= 16'hc5f;
assign q[10088]= 16'hd78;
assign q[10089]= 16'he57;
assign q[10090]= 16'hefd;
assign q[10091]= 16'hf6d;
assign q[10092]= 16'hfaa;
assign q[10093]= 16'hfbb;
assign q[10094]= 16'hfa7;
assign q[10095]= 16'hf77;
assign q[10096]= 16'hf33;
assign q[10097]= 16'hee6;
assign q[10098]= 16'he98;
assign q[10099]= 16'he53;
assign q[10100]= 16'he1e;
assign q[10101]= 16'he00;
assign q[10102]= 16'hdff;
assign q[10103]= 16'he1c;
assign q[10104]= 16'he58;
assign q[10105]= 16'heb4;
assign q[10106]= 16'hf2a;
assign q[10107]= 16'hfb5;
assign q[10108]= 16'h104f;
assign q[10109]= 16'h10ee;
assign q[10110]= 16'h1186;
assign q[10111]= 16'h120e;
assign q[10112]= 16'h1279;
assign q[10113]= 16'h12bb;
assign q[10114]= 16'h12c8;
assign q[10115]= 16'h1296;
assign q[10116]= 16'h121c;
assign q[10117]= 16'h1150;
assign q[10118]= 16'h102f;
assign q[10119]= 16'heb3;
assign q[10120]= 16'hcdb;
assign q[10121]= 16'haa9;
assign q[10122]= 16'h820;
assign q[10123]= 16'h547;
assign q[10124]= 16'h224;
assign q[10125]= 16'hfec4;
assign q[10126]= 16'hfb31;
assign q[10127]= 16'hf779;
assign q[10128]= 16'hf3aa;
assign q[10129]= 16'hefd4;
assign q[10130]= 16'hec07;
assign q[10131]= 16'he852;
assign q[10132]= 16'he4c4;
assign q[10133]= 16'he16d;
assign q[10134]= 16'hde5b;
assign q[10135]= 16'hdb99;
assign q[10136]= 16'hd935;
assign q[10137]= 16'hd736;
assign q[10138]= 16'hd5a7;
assign q[10139]= 16'hd48d;
assign q[10140]= 16'hd3ee;
assign q[10141]= 16'hd3cd;
assign q[10142]= 16'hd42b;
assign q[10143]= 16'hd50a;
assign q[10144]= 16'hd666;
assign q[10145]= 16'hd83e;
assign q[10146]= 16'hda8c;
assign q[10147]= 16'hdd4b;
assign q[10148]= 16'he073;
assign q[10149]= 16'he3fa;
assign q[10150]= 16'he7d8;
assign q[10151]= 16'hec00;
assign q[10152]= 16'hf066;
assign q[10153]= 16'hf4fc;
assign q[10154]= 16'hf9b3;
assign q[10155]= 16'hfe7c;
assign q[10156]= 16'h346;
assign q[10157]= 16'h801;
assign q[10158]= 16'hc9c;
assign q[10159]= 16'h1106;
assign q[10160]= 16'h152e;
assign q[10161]= 16'h1904;
assign q[10162]= 16'h1c78;
assign q[10163]= 16'h1f7c;
assign q[10164]= 16'h2205;
assign q[10165]= 16'h2407;
assign q[10166]= 16'h257a;
assign q[10167]= 16'h2659;
assign q[10168]= 16'h26a0;
assign q[10169]= 16'h264e;
assign q[10170]= 16'h2566;
assign q[10171]= 16'h23ed;
assign q[10172]= 16'h21ea;
assign q[10173]= 16'h1f68;
assign q[10174]= 16'h1c74;
assign q[10175]= 16'h191c;
assign q[10176]= 16'h156f;
assign q[10177]= 16'h1181;
assign q[10178]= 16'hd61;
assign q[10179]= 16'h924;
assign q[10180]= 16'h4d9;
assign q[10181]= 16'h93;
assign q[10182]= 16'hfc62;
assign q[10183]= 16'hf853;
assign q[10184]= 16'hf472;
assign q[10185]= 16'hf0cb;
assign q[10186]= 16'hed63;
assign q[10187]= 16'hea42;
assign q[10188]= 16'he768;
assign q[10189]= 16'he4d8;
assign q[10190]= 16'he28e;
assign q[10191]= 16'he088;
assign q[10192]= 16'hdebf;
assign q[10193]= 16'hdd2d;
assign q[10194]= 16'hdbcc;
assign q[10195]= 16'hda91;
assign q[10196]= 16'hd977;
assign q[10197]= 16'hd875;
assign q[10198]= 16'hd785;
assign q[10199]= 16'hd6a2;
assign q[10200]= 16'hd5c7;
assign q[10201]= 16'hd4f1;
assign q[10202]= 16'hd420;
assign q[10203]= 16'hd355;
assign q[10204]= 16'hd293;
assign q[10205]= 16'hd1de;
assign q[10206]= 16'hd13b;
assign q[10207]= 16'hd0b1;
assign q[10208]= 16'hd048;
assign q[10209]= 16'hd009;
assign q[10210]= 16'hcffb;
assign q[10211]= 16'hd026;
assign q[10212]= 16'hd093;
assign q[10213]= 16'hd148;
assign q[10214]= 16'hd24b;
assign q[10215]= 16'hd39f;
assign q[10216]= 16'hd547;
assign q[10217]= 16'hd743;
assign q[10218]= 16'hd993;
assign q[10219]= 16'hdc34;
assign q[10220]= 16'hdf1f;
assign q[10221]= 16'he24e;
assign q[10222]= 16'he5ba;
assign q[10223]= 16'he957;
assign q[10224]= 16'hed1b;
assign q[10225]= 16'hf0fa;
assign q[10226]= 16'hf4e7;
assign q[10227]= 16'hf8d5;
assign q[10228]= 16'hfcb8;
assign q[10229]= 16'h81;
assign q[10230]= 16'h425;
assign q[10231]= 16'h798;
assign q[10232]= 16'hacf;
assign q[10233]= 16'hdbf;
assign q[10234]= 16'h1060;
assign q[10235]= 16'h12aa;
assign q[10236]= 16'h1497;
assign q[10237]= 16'h1620;
assign q[10238]= 16'h1743;
assign q[10239]= 16'h17fd;
assign q[10240]= 16'h184d;
assign q[10241]= 16'h1832;
assign q[10242]= 16'h17ae;
assign q[10243]= 16'h16c4;
assign q[10244]= 16'h1576;
assign q[10245]= 16'h13c9;
assign q[10246]= 16'h11c3;
assign q[10247]= 16'hf69;
assign q[10248]= 16'hcc3;
assign q[10249]= 16'h9da;
assign q[10250]= 16'h6b4;
assign q[10251]= 16'h35d;
assign q[10252]= 16'hffde;
assign q[10253]= 16'hfc41;
assign q[10254]= 16'hf890;
assign q[10255]= 16'hf4d8;
assign q[10256]= 16'hf123;
assign q[10257]= 16'hed7e;
assign q[10258]= 16'he9f4;
assign q[10259]= 16'he68f;
assign q[10260]= 16'he35d;
assign q[10261]= 16'he066;
assign q[10262]= 16'hddb7;
assign q[10263]= 16'hdb57;
assign q[10264]= 16'hd950;
assign q[10265]= 16'hd7a9;
assign q[10266]= 16'hd66a;
assign q[10267]= 16'hd597;
assign q[10268]= 16'hd533;
assign q[10269]= 16'hd543;
assign q[10270]= 16'hd5c6;
assign q[10271]= 16'hd6bd;
assign q[10272]= 16'hd825;
assign q[10273]= 16'hd9fb;
assign q[10274]= 16'hdc3a;
assign q[10275]= 16'hdedc;
assign q[10276]= 16'he1d9;
assign q[10277]= 16'he529;
assign q[10278]= 16'he8c1;
assign q[10279]= 16'hec97;
assign q[10280]= 16'hf0a0;
assign q[10281]= 16'hf4d0;
assign q[10282]= 16'hf91a;
assign q[10283]= 16'hfd73;
assign q[10284]= 16'h1cb;
assign q[10285]= 16'h619;
assign q[10286]= 16'ha51;
assign q[10287]= 16'he65;
assign q[10288]= 16'h124b;
assign q[10289]= 16'h15fa;
assign q[10290]= 16'h1967;
assign q[10291]= 16'h1c8b;
assign q[10292]= 16'h1f5d;
assign q[10293]= 16'h21d8;
assign q[10294]= 16'h23f7;
assign q[10295]= 16'h25b6;
assign q[10296]= 16'h2713;
assign q[10297]= 16'h280c;
assign q[10298]= 16'h28a1;
assign q[10299]= 16'h28d2;
assign q[10300]= 16'h28a3;
assign q[10301]= 16'h2817;
assign q[10302]= 16'h2730;
assign q[10303]= 16'h25f5;
assign q[10304]= 16'h246c;
assign q[10305]= 16'h229a;
assign q[10306]= 16'h2087;
assign q[10307]= 16'h1e3b;
assign q[10308]= 16'h1bbe;
assign q[10309]= 16'h1918;
assign q[10310]= 16'h1653;
assign q[10311]= 16'h1376;
assign q[10312]= 16'h108d;
assign q[10313]= 16'hd9e;
assign q[10314]= 16'hab4;
assign q[10315]= 16'h7d8;
assign q[10316]= 16'h511;
assign q[10317]= 16'h269;
assign q[10318]= 16'hffe8;
assign q[10319]= 16'hfd93;
assign q[10320]= 16'hfb72;
assign q[10321]= 16'hf98c;
assign q[10322]= 16'hf7e5;
assign q[10323]= 16'hf682;
assign q[10324]= 16'hf568;
assign q[10325]= 16'hf497;
assign q[10326]= 16'hf413;
assign q[10327]= 16'hf3da;
assign q[10328]= 16'hf3ee;
assign q[10329]= 16'hf44b;
assign q[10330]= 16'hf4f0;
assign q[10331]= 16'hf5d7;
assign q[10332]= 16'hf6fc;
assign q[10333]= 16'hf85a;
assign q[10334]= 16'hf9e8;
assign q[10335]= 16'hfb9f;
assign q[10336]= 16'hfd77;
assign q[10337]= 16'hff68;
assign q[10338]= 16'h167;
assign q[10339]= 16'h36d;
assign q[10340]= 16'h570;
assign q[10341]= 16'h768;
assign q[10342]= 16'h94c;
assign q[10343]= 16'hb14;
assign q[10344]= 16'hcba;
assign q[10345]= 16'he37;
assign q[10346]= 16'hf87;
assign q[10347]= 16'h10a6;
assign q[10348]= 16'h1190;
assign q[10349]= 16'h1245;
assign q[10350]= 16'h12c3;
assign q[10351]= 16'h130b;
assign q[10352]= 16'h131d;
assign q[10353]= 16'h12fd;
assign q[10354]= 16'h12ab;
assign q[10355]= 16'h122c;
assign q[10356]= 16'h1183;
assign q[10357]= 16'h10b3;
assign q[10358]= 16'hfc0;
assign q[10359]= 16'head;
assign q[10360]= 16'hd7f;
assign q[10361]= 16'hc38;
assign q[10362]= 16'hadb;
assign q[10363]= 16'h96b;
assign q[10364]= 16'h7ea;
assign q[10365]= 16'h65a;
assign q[10366]= 16'h4bd;
assign q[10367]= 16'h315;
assign q[10368]= 16'h164;
assign q[10369]= 16'hffad;
assign q[10370]= 16'hfdf0;
assign q[10371]= 16'hfc30;
assign q[10372]= 16'hfa71;
assign q[10373]= 16'hf8b6;
assign q[10374]= 16'hf702;
assign q[10375]= 16'hf55b;
assign q[10376]= 16'hf3c4;
assign q[10377]= 16'hf244;
assign q[10378]= 16'hf0df;
assign q[10379]= 16'hef9c;
assign q[10380]= 16'hee80;
assign q[10381]= 16'hed90;
assign q[10382]= 16'hecd2;
assign q[10383]= 16'hec4a;
assign q[10384]= 16'hebfc;
assign q[10385]= 16'hebeb;
assign q[10386]= 16'hec19;
assign q[10387]= 16'hec86;
assign q[10388]= 16'hed33;
assign q[10389]= 16'hee1c;
assign q[10390]= 16'hef3f;
assign q[10391]= 16'hf098;
assign q[10392]= 16'hf220;
assign q[10393]= 16'hf3d2;
assign q[10394]= 16'hf5a5;
assign q[10395]= 16'hf791;
assign q[10396]= 16'hf98e;
assign q[10397]= 16'hfb93;
assign q[10398]= 16'hfd96;
assign q[10399]= 16'hff8e;
assign q[10400]= 16'h173;
assign q[10401]= 16'h33e;
assign q[10402]= 16'h4e6;
assign q[10403]= 16'h666;
assign q[10404]= 16'h7b7;
assign q[10405]= 16'h8d4;
assign q[10406]= 16'h9ba;
assign q[10407]= 16'ha65;
assign q[10408]= 16'had3;
assign q[10409]= 16'hb04;
assign q[10410]= 16'haf6;
assign q[10411]= 16'haa9;
assign q[10412]= 16'ha1e;
assign q[10413]= 16'h956;
assign q[10414]= 16'h853;
assign q[10415]= 16'h718;
assign q[10416]= 16'h5a7;
assign q[10417]= 16'h403;
assign q[10418]= 16'h232;
assign q[10419]= 16'h38;
assign q[10420]= 16'hfe1b;
assign q[10421]= 16'hfbe0;
assign q[10422]= 16'hf990;
assign q[10423]= 16'hf733;
assign q[10424]= 16'hf4d4;
assign q[10425]= 16'hf27c;
assign q[10426]= 16'hf037;
assign q[10427]= 16'hee11;
assign q[10428]= 16'hec18;
assign q[10429]= 16'hea58;
assign q[10430]= 16'he8df;
assign q[10431]= 16'he7ba;
assign q[10432]= 16'he6f5;
assign q[10433]= 16'he69b;
assign q[10434]= 16'he6b6;
assign q[10435]= 16'he74d;
assign q[10436]= 16'he866;
assign q[10437]= 16'hea03;
assign q[10438]= 16'hec23;
assign q[10439]= 16'heec3;
assign q[10440]= 16'hf1db;
assign q[10441]= 16'hf560;
assign q[10442]= 16'hf945;
assign q[10443]= 16'hfd77;
assign q[10444]= 16'h1e2;
assign q[10445]= 16'h672;
assign q[10446]= 16'hb0c;
assign q[10447]= 16'hf98;
assign q[10448]= 16'h13fb;
assign q[10449]= 16'h181c;
assign q[10450]= 16'h1be1;
assign q[10451]= 16'h1f34;
assign q[10452]= 16'h2201;
assign q[10453]= 16'h2435;
assign q[10454]= 16'h25c4;
assign q[10455]= 16'h26a4;
assign q[10456]= 16'h26d1;
assign q[10457]= 16'h264a;
assign q[10458]= 16'h2514;
assign q[10459]= 16'h2338;
assign q[10460]= 16'h20c5;
assign q[10461]= 16'h1dcd;
assign q[10462]= 16'h1a64;
assign q[10463]= 16'h16a4;
assign q[10464]= 16'h12a6;
assign q[10465]= 16'he86;
assign q[10466]= 16'ha60;
assign q[10467]= 16'h650;
assign q[10468]= 16'h26f;
assign q[10469]= 16'hfed9;
assign q[10470]= 16'hfb9f;
assign q[10471]= 16'hf8d6;
assign q[10472]= 16'hf68d;
assign q[10473]= 16'hf4cd;
assign q[10474]= 16'hf39f;
assign q[10475]= 16'hf303;
assign q[10476]= 16'hf2f8;
assign q[10477]= 16'hf379;
assign q[10478]= 16'hf47b;
assign q[10479]= 16'hf5f2;
assign q[10480]= 16'hf7ce;
assign q[10481]= 16'hf9ff;
assign q[10482]= 16'hfc71;
assign q[10483]= 16'hff12;
assign q[10484]= 16'h1cb;
assign q[10485]= 16'h48c;
assign q[10486]= 16'h742;
assign q[10487]= 16'h9db;
assign q[10488]= 16'hc48;
assign q[10489]= 16'he7e;
assign q[10490]= 16'h1070;
assign q[10491]= 16'h1218;
assign q[10492]= 16'h136f;
assign q[10493]= 16'h1474;
assign q[10494]= 16'h1525;
assign q[10495]= 16'h1585;
assign q[10496]= 16'h1597;
assign q[10497]= 16'h1562;
assign q[10498]= 16'h14ec;
assign q[10499]= 16'h143f;
assign q[10500]= 16'h1363;
assign q[10501]= 16'h1263;
assign q[10502]= 16'h1148;
assign q[10503]= 16'h101f;
assign q[10504]= 16'hef1;
assign q[10505]= 16'hdc8;
assign q[10506]= 16'hcae;
assign q[10507]= 16'hbab;
assign q[10508]= 16'hac9;
assign q[10509]= 16'ha0e;
assign q[10510]= 16'h980;
assign q[10511]= 16'h924;
assign q[10512]= 16'h900;
assign q[10513]= 16'h915;
assign q[10514]= 16'h966;
assign q[10515]= 16'h9f3;
assign q[10516]= 16'habc;
assign q[10517]= 16'hbbe;
assign q[10518]= 16'hcf8;
assign q[10519]= 16'he64;
assign q[10520]= 16'hffd;
assign q[10521]= 16'h11be;
assign q[10522]= 16'h13a0;
assign q[10523]= 16'h159a;
assign q[10524]= 16'h17a4;
assign q[10525]= 16'h19b5;
assign q[10526]= 16'h1bc4;
assign q[10527]= 16'h1dc7;
assign q[10528]= 16'h1fb5;
assign q[10529]= 16'h2186;
assign q[10530]= 16'h2330;
assign q[10531]= 16'h24ac;
assign q[10532]= 16'h25f3;
assign q[10533]= 16'h26ff;
assign q[10534]= 16'h27cb;
assign q[10535]= 16'h2854;
assign q[10536]= 16'h2898;
assign q[10537]= 16'h2895;
assign q[10538]= 16'h284d;
assign q[10539]= 16'h27c1;
assign q[10540]= 16'h26f4;
assign q[10541]= 16'h25ea;
assign q[10542]= 16'h24a9;
assign q[10543]= 16'h2336;
assign q[10544]= 16'h2197;
assign q[10545]= 16'h1fd5;
assign q[10546]= 16'h1df6;
assign q[10547]= 16'h1c02;
assign q[10548]= 16'h1a02;
assign q[10549]= 16'h17fc;
assign q[10550]= 16'h15fa;
assign q[10551]= 16'h1401;
assign q[10552]= 16'h121b;
assign q[10553]= 16'h104e;
assign q[10554]= 16'hea1;
assign q[10555]= 16'hd19;
assign q[10556]= 16'hbbe;
assign q[10557]= 16'ha94;
assign q[10558]= 16'h99f;
assign q[10559]= 16'h8e5;
assign q[10560]= 16'h868;
assign q[10561]= 16'h82a;
assign q[10562]= 16'h82d;
assign q[10563]= 16'h870;
assign q[10564]= 16'h8f3;
assign q[10565]= 16'h9b3;
assign q[10566]= 16'haaa;
assign q[10567]= 16'hbd4;
assign q[10568]= 16'hd27;
assign q[10569]= 16'he9a;
assign q[10570]= 16'h1021;
assign q[10571]= 16'h11b0;
assign q[10572]= 16'h1338;
assign q[10573]= 16'h14aa;
assign q[10574]= 16'h15f4;
assign q[10575]= 16'h1707;
assign q[10576]= 16'h17d3;
assign q[10577]= 16'h1846;
assign q[10578]= 16'h1853;
assign q[10579]= 16'h17ee;
assign q[10580]= 16'h170c;
assign q[10581]= 16'h15a6;
assign q[10582]= 16'h13b9;
assign q[10583]= 16'h1144;
assign q[10584]= 16'he4c;
assign q[10585]= 16'hada;
assign q[10586]= 16'h6fa;
assign q[10587]= 16'h2bd;
assign q[10588]= 16'hfe3a;
assign q[10589]= 16'hf986;
assign q[10590]= 16'hf4be;
assign q[10591]= 16'heffe;
assign q[10592]= 16'heb64;
assign q[10593]= 16'he70e;
assign q[10594]= 16'he31b;
assign q[10595]= 16'hdfa5;
assign q[10596]= 16'hdcc5;
assign q[10597]= 16'hda91;
assign q[10598]= 16'hd918;
assign q[10599]= 16'hd865;
assign q[10600]= 16'hd87f;
assign q[10601]= 16'hd964;
assign q[10602]= 16'hdb0c;
assign q[10603]= 16'hdd6b;
assign q[10604]= 16'he06d;
assign q[10605]= 16'he3f9;
assign q[10606]= 16'he7f2;
assign q[10607]= 16'hec38;
assign q[10608]= 16'hf0a5;
assign q[10609]= 16'hf515;
assign q[10610]= 16'hf963;
assign q[10611]= 16'hfd6a;
assign q[10612]= 16'h107;
assign q[10613]= 16'h41d;
assign q[10614]= 16'h690;
assign q[10615]= 16'h84d;
assign q[10616]= 16'h944;
assign q[10617]= 16'h96d;
assign q[10618]= 16'h8c6;
assign q[10619]= 16'h756;
assign q[10620]= 16'h528;
assign q[10621]= 16'h24f;
assign q[10622]= 16'hfee4;
assign q[10623]= 16'hfb03;
assign q[10624]= 16'hf6cb;
assign q[10625]= 16'hf262;
assign q[10626]= 16'hedea;
assign q[10627]= 16'he989;
assign q[10628]= 16'he562;
assign q[10629]= 16'he198;
assign q[10630]= 16'hde48;
assign q[10631]= 16'hdb8d;
assign q[10632]= 16'hd97d;
assign q[10633]= 16'hd828;
assign q[10634]= 16'hd799;
assign q[10635]= 16'hd7d5;
assign q[10636]= 16'hd8db;
assign q[10637]= 16'hdaa5;
assign q[10638]= 16'hdd28;
assign q[10639]= 16'he054;
assign q[10640]= 16'he415;
assign q[10641]= 16'he857;
assign q[10642]= 16'hecff;
assign q[10643]= 16'hf1f5;
assign q[10644]= 16'hf71e;
assign q[10645]= 16'hfc61;
assign q[10646]= 16'h1a3;
assign q[10647]= 16'h6cf;
assign q[10648]= 16'hbd0;
assign q[10649]= 16'h1092;
assign q[10650]= 16'h1507;
assign q[10651]= 16'h1921;
assign q[10652]= 16'h1cd6;
assign q[10653]= 16'h201f;
assign q[10654]= 16'h22f9;
assign q[10655]= 16'h2562;
assign q[10656]= 16'h2759;
assign q[10657]= 16'h28e1;
assign q[10658]= 16'h29ff;
assign q[10659]= 16'h2ab6;
assign q[10660]= 16'h2b0e;
assign q[10661]= 16'h2b0c;
assign q[10662]= 16'h2ab8;
assign q[10663]= 16'h2a1a;
assign q[10664]= 16'h293a;
assign q[10665]= 16'h281e;
assign q[10666]= 16'h26d0;
assign q[10667]= 16'h2556;
assign q[10668]= 16'h23ba;
assign q[10669]= 16'h2203;
assign q[10670]= 16'h2039;
assign q[10671]= 16'h1e64;
assign q[10672]= 16'h1c8d;
assign q[10673]= 16'h1abc;
assign q[10674]= 16'h18f9;
assign q[10675]= 16'h174a;
assign q[10676]= 16'h15b8;
assign q[10677]= 16'h1449;
assign q[10678]= 16'h1302;
assign q[10679]= 16'h11e8;
assign q[10680]= 16'h10fd;
assign q[10681]= 16'h1043;
assign q[10682]= 16'hfbb;
assign q[10683]= 16'hf62;
assign q[10684]= 16'hf34;
assign q[10685]= 16'hf2c;
assign q[10686]= 16'hf42;
assign q[10687]= 16'hf6f;
assign q[10688]= 16'hfa8;
assign q[10689]= 16'hfe1;
assign q[10690]= 16'h1011;
assign q[10691]= 16'h102b;
assign q[10692]= 16'h1025;
assign q[10693]= 16'hff4;
assign q[10694]= 16'hf8f;
assign q[10695]= 16'hef0;
assign q[10696]= 16'he12;
assign q[10697]= 16'hcf2;
assign q[10698]= 16'hb91;
assign q[10699]= 16'h9f2;
assign q[10700]= 16'h81b;
assign q[10701]= 16'h615;
assign q[10702]= 16'h3eb;
assign q[10703]= 16'h1aa;
assign q[10704]= 16'hff62;
assign q[10705]= 16'hfd22;
assign q[10706]= 16'hfafb;
assign q[10707]= 16'hf8ff;
assign q[10708]= 16'hf73c;
assign q[10709]= 16'hf5c3;
assign q[10710]= 16'hf49f;
assign q[10711]= 16'hf3db;
assign q[10712]= 16'hf37f;
assign q[10713]= 16'hf38e;
assign q[10714]= 16'hf408;
assign q[10715]= 16'hf4eb;
assign q[10716]= 16'hf630;
assign q[10717]= 16'hf7cb;
assign q[10718]= 16'hf9b0;
assign q[10719]= 16'hfbcf;
assign q[10720]= 16'hfe15;
assign q[10721]= 16'h6d;
assign q[10722]= 16'h2c4;
assign q[10723]= 16'h505;
assign q[10724]= 16'h71b;
assign q[10725]= 16'h8f4;
assign q[10726]= 16'ha7f;
assign q[10727]= 16'hbad;
assign q[10728]= 16'hc74;
assign q[10729]= 16'hccd;
assign q[10730]= 16'hcb3;
assign q[10731]= 16'hc28;
assign q[10732]= 16'hb2f;
assign q[10733]= 16'h9d1;
assign q[10734]= 16'h819;
assign q[10735]= 16'h617;
assign q[10736]= 16'h3db;
assign q[10737]= 16'h179;
assign q[10738]= 16'hff06;
assign q[10739]= 16'hfc96;
assign q[10740]= 16'hfa3e;
assign q[10741]= 16'hf813;
assign q[10742]= 16'hf626;
assign q[10743]= 16'hf48a;
assign q[10744]= 16'hf34a;
assign q[10745]= 16'hf274;
assign q[10746]= 16'hf20d;
assign q[10747]= 16'hf21a;
assign q[10748]= 16'hf29c;
assign q[10749]= 16'hf38f;
assign q[10750]= 16'hf4ef;
assign q[10751]= 16'hf6b2;
assign q[10752]= 16'hf8cd;
assign q[10753]= 16'hfb33;
assign q[10754]= 16'hfdd5;
assign q[10755]= 16'ha2;
assign q[10756]= 16'h38d;
assign q[10757]= 16'h686;
assign q[10758]= 16'h97d;
assign q[10759]= 16'hc67;
assign q[10760]= 16'hf36;
assign q[10761]= 16'h11e2;
assign q[10762]= 16'h1464;
assign q[10763]= 16'h16b7;
assign q[10764]= 16'h18d7;
assign q[10765]= 16'h1ac5;
assign q[10766]= 16'h1c83;
assign q[10767]= 16'h1e13;
assign q[10768]= 16'h1f79;
assign q[10769]= 16'h20bd;
assign q[10770]= 16'h21e2;
assign q[10771]= 16'h22ef;
assign q[10772]= 16'h23e9;
assign q[10773]= 16'h24d3;
assign q[10774]= 16'h25b0;
assign q[10775]= 16'h2680;
assign q[10776]= 16'h2742;
assign q[10777]= 16'h27f2;
assign q[10778]= 16'h288b;
assign q[10779]= 16'h2905;
assign q[10780]= 16'h2955;
assign q[10781]= 16'h2971;
assign q[10782]= 16'h294d;
assign q[10783]= 16'h28db;
assign q[10784]= 16'h280f;
assign q[10785]= 16'h26dc;
assign q[10786]= 16'h2539;
assign q[10787]= 16'h231c;
assign q[10788]= 16'h2081;
assign q[10789]= 16'h1d63;
assign q[10790]= 16'h19c5;
assign q[10791]= 16'h15ab;
assign q[10792]= 16'h111f;
assign q[10793]= 16'hc30;
assign q[10794]= 16'h6ef;
assign q[10795]= 16'h173;
assign q[10796]= 16'hfbd6;
assign q[10797]= 16'hf635;
assign q[10798]= 16'hf0af;
assign q[10799]= 16'heb65;
assign q[10800]= 16'he678;
assign q[10801]= 16'he209;
assign q[10802]= 16'hde36;
assign q[10803]= 16'hdb1d;
assign q[10804]= 16'hd8d5;
assign q[10805]= 16'hd771;
assign q[10806]= 16'hd701;
assign q[10807]= 16'hd78c;
assign q[10808]= 16'hd912;
assign q[10809]= 16'hdb8f;
assign q[10810]= 16'hdef5;
assign q[10811]= 16'he330;
assign q[10812]= 16'he825;
assign q[10813]= 16'hedb5;
assign q[10814]= 16'hf3b9;
assign q[10815]= 16'hfa09;
assign q[10816]= 16'h77;
assign q[10817]= 16'h6d7;
assign q[10818]= 16'hcf9;
assign q[10819]= 16'h12b2;
assign q[10820]= 16'h17d7;
assign q[10821]= 16'h1c42;
assign q[10822]= 16'h1fd2;
assign q[10823]= 16'h226b;
assign q[10824]= 16'h23f9;
assign q[10825]= 16'h2471;
assign q[10826]= 16'h23ce;
assign q[10827]= 16'h2213;
assign q[10828]= 16'h1f4d;
assign q[10829]= 16'h1b8d;
assign q[10830]= 16'h16ee;
assign q[10831]= 16'h118f;
assign q[10832]= 16'hb95;
assign q[10833]= 16'h527;
assign q[10834]= 16'hfe72;
assign q[10835]= 16'hf79c;
assign q[10836]= 16'hf0d3;
assign q[10837]= 16'hea3e;
assign q[10838]= 16'he402;
assign q[10839]= 16'hde41;
assign q[10840]= 16'hd914;
assign q[10841]= 16'hd493;
assign q[10842]= 16'hd0cc;
assign q[10843]= 16'hcdc7;
assign q[10844]= 16'hcb86;
assign q[10845]= 16'hca04;
assign q[10846]= 16'hc936;
assign q[10847]= 16'hc90d;
assign q[10848]= 16'hc974;
assign q[10849]= 16'hca52;
assign q[10850]= 16'hcb8e;
assign q[10851]= 16'hcd0d;
assign q[10852]= 16'hceb3;
assign q[10853]= 16'hd066;
assign q[10854]= 16'hd20e;
assign q[10855]= 16'hd395;
assign q[10856]= 16'hd4e9;
assign q[10857]= 16'hd5fe;
assign q[10858]= 16'hd6cb;
assign q[10859]= 16'hd74a;
assign q[10860]= 16'hd77d;
assign q[10861]= 16'hd768;
assign q[10862]= 16'hd714;
assign q[10863]= 16'hd68c;
assign q[10864]= 16'hd5e0;
assign q[10865]= 16'hd51f;
assign q[10866]= 16'hd45b;
assign q[10867]= 16'hd3a5;
assign q[10868]= 16'hd30e;
assign q[10869]= 16'hd2a5;
assign q[10870]= 16'hd278;
assign q[10871]= 16'hd291;
assign q[10872]= 16'hd2f7;
assign q[10873]= 16'hd3af;
assign q[10874]= 16'hd4b8;
assign q[10875]= 16'hd611;
assign q[10876]= 16'hd7b3;
assign q[10877]= 16'hd996;
assign q[10878]= 16'hdbae;
assign q[10879]= 16'hddef;
assign q[10880]= 16'he04b;
assign q[10881]= 16'he2b1;
assign q[10882]= 16'he514;
assign q[10883]= 16'he766;
assign q[10884]= 16'he999;
assign q[10885]= 16'heba2;
assign q[10886]= 16'hed78;
assign q[10887]= 16'hef13;
assign q[10888]= 16'hf06f;
assign q[10889]= 16'hf189;
assign q[10890]= 16'hf263;
assign q[10891]= 16'hf2fe;
assign q[10892]= 16'hf360;
assign q[10893]= 16'hf38d;
assign q[10894]= 16'hf38f;
assign q[10895]= 16'hf36d;
assign q[10896]= 16'hf330;
assign q[10897]= 16'hf2e1;
assign q[10898]= 16'hf287;
assign q[10899]= 16'hf22b;
assign q[10900]= 16'hf1d4;
assign q[10901]= 16'hf185;
assign q[10902]= 16'hf143;
assign q[10903]= 16'hf111;
assign q[10904]= 16'hf0f0;
assign q[10905]= 16'hf0df;
assign q[10906]= 16'hf0dc;
assign q[10907]= 16'hf0e7;
assign q[10908]= 16'hf0fa;
assign q[10909]= 16'hf114;
assign q[10910]= 16'hf130;
assign q[10911]= 16'hf14b;
assign q[10912]= 16'hf162;
assign q[10913]= 16'hf171;
assign q[10914]= 16'hf178;
assign q[10915]= 16'hf175;
assign q[10916]= 16'hf168;
assign q[10917]= 16'hf151;
assign q[10918]= 16'hf131;
assign q[10919]= 16'hf10a;
assign q[10920]= 16'hf0df;
assign q[10921]= 16'hf0b3;
assign q[10922]= 16'hf088;
assign q[10923]= 16'hf062;
assign q[10924]= 16'hf043;
assign q[10925]= 16'hf02e;
assign q[10926]= 16'hf026;
assign q[10927]= 16'hf02c;
assign q[10928]= 16'hf041;
assign q[10929]= 16'hf066;
assign q[10930]= 16'hf09c;
assign q[10931]= 16'hf0e2;
assign q[10932]= 16'hf139;
assign q[10933]= 16'hf1a0;
assign q[10934]= 16'hf218;
assign q[10935]= 16'hf2a0;
assign q[10936]= 16'hf338;
assign q[10937]= 16'hf3e2;
assign q[10938]= 16'hf49f;
assign q[10939]= 16'hf570;
assign q[10940]= 16'hf65a;
assign q[10941]= 16'hf75d;
assign q[10942]= 16'hf87f;
assign q[10943]= 16'hf9c1;
assign q[10944]= 16'hfb29;
assign q[10945]= 16'hfcb9;
assign q[10946]= 16'hfe74;
assign q[10947]= 16'h5c;
assign q[10948]= 16'h272;
assign q[10949]= 16'h4b7;
assign q[10950]= 16'h727;
assign q[10951]= 16'h9c1;
assign q[10952]= 16'hc7f;
assign q[10953]= 16'hf5a;
assign q[10954]= 16'h124a;
assign q[10955]= 16'h1544;
assign q[10956]= 16'h183d;
assign q[10957]= 16'h1b29;
assign q[10958]= 16'h1dfb;
assign q[10959]= 16'h20a4;
assign q[10960]= 16'h2317;
assign q[10961]= 16'h2547;
assign q[10962]= 16'h2728;
assign q[10963]= 16'h28b1;
assign q[10964]= 16'h29d7;
assign q[10965]= 16'h2a95;
assign q[10966]= 16'h2ae8;
assign q[10967]= 16'h2ace;
assign q[10968]= 16'h2a4a;
assign q[10969]= 16'h2961;
assign q[10970]= 16'h281b;
assign q[10971]= 16'h2683;
assign q[10972]= 16'h24a6;
assign q[10973]= 16'h2295;
assign q[10974]= 16'h2060;
assign q[10975]= 16'h1e1a;
assign q[10976]= 16'h1bd5;
assign q[10977]= 16'h19a5;
assign q[10978]= 16'h179c;
assign q[10979]= 16'h15ca;
assign q[10980]= 16'h1440;
assign q[10981]= 16'h1309;
assign q[10982]= 16'h1230;
assign q[10983]= 16'h11bc;
assign q[10984]= 16'h11b1;
assign q[10985]= 16'h120e;
assign q[10986]= 16'h12d0;
assign q[10987]= 16'h13f0;
assign q[10988]= 16'h1565;
assign q[10989]= 16'h1720;
assign q[10990]= 16'h1912;
assign q[10991]= 16'h1b2a;
assign q[10992]= 16'h1d53;
assign q[10993]= 16'h1f7a;
assign q[10994]= 16'h218b;
assign q[10995]= 16'h2370;
assign q[10996]= 16'h2516;
assign q[10997]= 16'h266c;
assign q[10998]= 16'h2761;
assign q[10999]= 16'h27e9;
assign q[11000]= 16'h27f7;
assign q[11001]= 16'h2785;
assign q[11002]= 16'h268f;
assign q[11003]= 16'h2514;
assign q[11004]= 16'h2316;
assign q[11005]= 16'h209c;
assign q[11006]= 16'h1dae;
assign q[11007]= 16'h1a59;
assign q[11008]= 16'h16ac;
assign q[11009]= 16'h12b6;
assign q[11010]= 16'he8b;
assign q[11011]= 16'ha3e;
assign q[11012]= 16'h5e2;
assign q[11013]= 16'h18c;
assign q[11014]= 16'hfd52;
assign q[11015]= 16'hf943;
assign q[11016]= 16'hf574;
assign q[11017]= 16'hf1f4;
assign q[11018]= 16'heed2;
assign q[11019]= 16'hec19;
assign q[11020]= 16'he9d5;
assign q[11021]= 16'he80d;
assign q[11022]= 16'he6c4;
assign q[11023]= 16'he5ff;
assign q[11024]= 16'he5bc;
assign q[11025]= 16'he5fb;
assign q[11026]= 16'he6b6;
assign q[11027]= 16'he7e7;
assign q[11028]= 16'he988;
assign q[11029]= 16'heb8e;
assign q[11030]= 16'hedf0;
assign q[11031]= 16'hf0a3;
assign q[11032]= 16'hf39c;
assign q[11033]= 16'hf6cf;
assign q[11034]= 16'hfa30;
assign q[11035]= 16'hfdb4;
assign q[11036]= 16'h14e;
assign q[11037]= 16'h4f6;
assign q[11038]= 16'h89f;
assign q[11039]= 16'hc40;
assign q[11040]= 16'hfcf;
assign q[11041]= 16'h1343;
assign q[11042]= 16'h1695;
assign q[11043]= 16'h19bb;
assign q[11044]= 16'h1caf;
assign q[11045]= 16'h1f69;
assign q[11046]= 16'h21e2;
assign q[11047]= 16'h2414;
assign q[11048]= 16'h25f8;
assign q[11049]= 16'h278a;
assign q[11050]= 16'h28c2;
assign q[11051]= 16'h299d;
assign q[11052]= 16'h2a15;
assign q[11053]= 16'h2a27;
assign q[11054]= 16'h29cf;
assign q[11055]= 16'h290b;
assign q[11056]= 16'h27db;
assign q[11057]= 16'h263d;
assign q[11058]= 16'h2434;
assign q[11059]= 16'h21c3;
assign q[11060]= 16'h1eed;
assign q[11061]= 16'h1bb9;
assign q[11062]= 16'h182e;
assign q[11063]= 16'h1456;
assign q[11064]= 16'h103c;
assign q[11065]= 16'hbec;
assign q[11066]= 16'h774;
assign q[11067]= 16'h2e1;
assign q[11068]= 16'hfe46;
assign q[11069]= 16'hf9af;
assign q[11070]= 16'hf52d;
assign q[11071]= 16'hf0d0;
assign q[11072]= 16'heca8;
assign q[11073]= 16'he8c2;
assign q[11074]= 16'he52c;
assign q[11075]= 16'he1f1;
assign q[11076]= 16'hdf1b;
assign q[11077]= 16'hdcb1;
assign q[11078]= 16'hdab8;
assign q[11079]= 16'hd935;
assign q[11080]= 16'hd827;
assign q[11081]= 16'hd78d;
assign q[11082]= 16'hd763;
assign q[11083]= 16'hd7a4;
assign q[11084]= 16'hd849;
assign q[11085]= 16'hd947;
assign q[11086]= 16'hda97;
assign q[11087]= 16'hdc2b;
assign q[11088]= 16'hddfa;
assign q[11089]= 16'hdff8;
assign q[11090]= 16'he219;
assign q[11091]= 16'he453;
assign q[11092]= 16'he69d;
assign q[11093]= 16'he8ed;
assign q[11094]= 16'heb3c;
assign q[11095]= 16'hed84;
assign q[11096]= 16'hefc1;
assign q[11097]= 16'hf1ef;
assign q[11098]= 16'hf40c;
assign q[11099]= 16'hf619;
assign q[11100]= 16'hf815;
assign q[11101]= 16'hfa03;
assign q[11102]= 16'hfbe5;
assign q[11103]= 16'hfdbd;
assign q[11104]= 16'hff8f;
assign q[11105]= 16'h15d;
assign q[11106]= 16'h32c;
assign q[11107]= 16'h4fe;
assign q[11108]= 16'h6d5;
assign q[11109]= 16'h8b2;
assign q[11110]= 16'ha97;
assign q[11111]= 16'hc83;
assign q[11112]= 16'he76;
assign q[11113]= 16'h106f;
assign q[11114]= 16'h126c;
assign q[11115]= 16'h1469;
assign q[11116]= 16'h1665;
assign q[11117]= 16'h185b;
assign q[11118]= 16'h1a48;
assign q[11119]= 16'h1c28;
assign q[11120]= 16'h1df7;
assign q[11121]= 16'h1fb2;
assign q[11122]= 16'h2154;
assign q[11123]= 16'h22d9;
assign q[11124]= 16'h243e;
assign q[11125]= 16'h257f;
assign q[11126]= 16'h2698;
assign q[11127]= 16'h2786;
assign q[11128]= 16'h2844;
assign q[11129]= 16'h28cf;
assign q[11130]= 16'h2923;
assign q[11131]= 16'h293d;
assign q[11132]= 16'h2918;
assign q[11133]= 16'h28b1;
assign q[11134]= 16'h2804;
assign q[11135]= 16'h270f;
assign q[11136]= 16'h25ce;
assign q[11137]= 16'h2440;
assign q[11138]= 16'h2265;
assign q[11139]= 16'h203d;
assign q[11140]= 16'h1dc9;
assign q[11141]= 16'h1b0e;
assign q[11142]= 16'h1811;
assign q[11143]= 16'h14da;
assign q[11144]= 16'h1172;
assign q[11145]= 16'hde5;
assign q[11146]= 16'ha41;
assign q[11147]= 16'h696;
assign q[11148]= 16'h2f5;
assign q[11149]= 16'hff71;
assign q[11150]= 16'hfc1c;
assign q[11151]= 16'hf90b;
assign q[11152]= 16'hf652;
assign q[11153]= 16'hf402;
assign q[11154]= 16'hf22e;
assign q[11155]= 16'hf0e5;
assign q[11156]= 16'hf032;
assign q[11157]= 16'hf020;
assign q[11158]= 16'hf0b3;
assign q[11159]= 16'hf1ed;
assign q[11160]= 16'hf3ca;
assign q[11161]= 16'hf642;
assign q[11162]= 16'hf948;
assign q[11163]= 16'hfccc;
assign q[11164]= 16'hb7;
assign q[11165]= 16'h4f2;
assign q[11166]= 16'h960;
assign q[11167]= 16'hde4;
assign q[11168]= 16'h125c;
assign q[11169]= 16'h16aa;
assign q[11170]= 16'h1aad;
assign q[11171]= 16'h1e48;
assign q[11172]= 16'h215f;
assign q[11173]= 16'h23db;
assign q[11174]= 16'h25a8;
assign q[11175]= 16'h26b7;
assign q[11176]= 16'h2700;
assign q[11177]= 16'h2681;
assign q[11178]= 16'h253c;
assign q[11179]= 16'h233c;
assign q[11180]= 16'h2092;
assign q[11181]= 16'h1d51;
assign q[11182]= 16'h1996;
assign q[11183]= 16'h157d;
assign q[11184]= 16'h112b;
assign q[11185]= 16'hcc1;
assign q[11186]= 16'h865;
assign q[11187]= 16'h43d;
assign q[11188]= 16'h6a;
assign q[11189]= 16'hfd0e;
assign q[11190]= 16'hfa44;
assign q[11191]= 16'hf825;
assign q[11192]= 16'hf6c3;
assign q[11193]= 16'hf62b;
assign q[11194]= 16'hf663;
assign q[11195]= 16'hf76a;
assign q[11196]= 16'hf939;
assign q[11197]= 16'hfbc1;
assign q[11198]= 16'hfef0;
assign q[11199]= 16'h2aa;
assign q[11200]= 16'h6d7;
assign q[11201]= 16'hb53;
assign q[11202]= 16'hffc;
assign q[11203]= 16'h14af;
assign q[11204]= 16'h1949;
assign q[11205]= 16'h1da7;
assign q[11206]= 16'h21aa;
assign q[11207]= 16'h2536;
assign q[11208]= 16'h2833;
assign q[11209]= 16'h2a8f;
assign q[11210]= 16'h2c3d;
assign q[11211]= 16'h2d34;
assign q[11212]= 16'h2d75;
assign q[11213]= 16'h2d02;
assign q[11214]= 16'h2be7;
assign q[11215]= 16'h2a31;
assign q[11216]= 16'h27f3;
assign q[11217]= 16'h2542;
assign q[11218]= 16'h2239;
assign q[11219]= 16'h1eef;
assign q[11220]= 16'h1b7f;
assign q[11221]= 16'h1802;
assign q[11222]= 16'h148f;
assign q[11223]= 16'h113c;
assign q[11224]= 16'he19;
assign q[11225]= 16'hb36;
assign q[11226]= 16'h89b;
assign q[11227]= 16'h64e;
assign q[11228]= 16'h44f;
assign q[11229]= 16'h29b;
assign q[11230]= 16'h129;
assign q[11231]= 16'hfff1;
assign q[11232]= 16'hfee1;
assign q[11233]= 16'hfdeb;
assign q[11234]= 16'hfcff;
assign q[11235]= 16'hfc0a;
assign q[11236]= 16'hfafe;
assign q[11237]= 16'hf9ca;
assign q[11238]= 16'hf863;
assign q[11239]= 16'hf6be;
assign q[11240]= 16'hf4d6;
assign q[11241]= 16'hf2aa;
assign q[11242]= 16'hf03b;
assign q[11243]= 16'hed90;
assign q[11244]= 16'heab4;
assign q[11245]= 16'he7b5;
assign q[11246]= 16'he4a4;
assign q[11247]= 16'he196;
assign q[11248]= 16'hde9f;
assign q[11249]= 16'hdbd7;
assign q[11250]= 16'hd953;
assign q[11251]= 16'hd729;
assign q[11252]= 16'hd56b;
assign q[11253]= 16'hd428;
assign q[11254]= 16'hd36d;
assign q[11255]= 16'hd341;
assign q[11256]= 16'hd3a7;
assign q[11257]= 16'hd49b;
assign q[11258]= 16'hd616;
assign q[11259]= 16'hd80a;
assign q[11260]= 16'hda66;
assign q[11261]= 16'hdd12;
assign q[11262]= 16'hdff5;
assign q[11263]= 16'he2f2;
assign q[11264]= 16'he5ec;
assign q[11265]= 16'he8c4;
assign q[11266]= 16'heb5c;
assign q[11267]= 16'hed9a;
assign q[11268]= 16'hef64;
assign q[11269]= 16'hf0a6;
assign q[11270]= 16'hf152;
assign q[11271]= 16'hf15d;
assign q[11272]= 16'hf0c6;
assign q[11273]= 16'hef8f;
assign q[11274]= 16'hedc4;
assign q[11275]= 16'heb75;
assign q[11276]= 16'he8ba;
assign q[11277]= 16'he5af;
assign q[11278]= 16'he276;
assign q[11279]= 16'hdf31;
assign q[11280]= 16'hdc07;
assign q[11281]= 16'hd920;
assign q[11282]= 16'hd6a0;
assign q[11283]= 16'hd4ac;
assign q[11284]= 16'hd362;
assign q[11285]= 16'hd2df;
assign q[11286]= 16'hd336;
assign q[11287]= 16'hd475;
assign q[11288]= 16'hd6a2;
assign q[11289]= 16'hd9ba;
assign q[11290]= 16'hddb2;
assign q[11291]= 16'he279;
assign q[11292]= 16'he7f2;
assign q[11293]= 16'hedfe;
assign q[11294]= 16'hf473;
assign q[11295]= 16'hfb27;
assign q[11296]= 16'h1e9;
assign q[11297]= 16'h88a;
assign q[11298]= 16'hed8;
assign q[11299]= 16'h14a5;
assign q[11300]= 16'h19c4;
assign q[11301]= 16'h1e0e;
assign q[11302]= 16'h2162;
assign q[11303]= 16'h23a7;
assign q[11304]= 16'h24cb;
assign q[11305]= 16'h24c6;
assign q[11306]= 16'h2397;
assign q[11307]= 16'h2149;
assign q[11308]= 16'h1ded;
assign q[11309]= 16'h199d;
assign q[11310]= 16'h147c;
assign q[11311]= 16'heaf;
assign q[11312]= 16'h864;
assign q[11313]= 16'h1c9;
assign q[11314]= 16'hfb0f;
assign q[11315]= 16'hf465;
assign q[11316]= 16'hedfb;
assign q[11317]= 16'he7fb;
assign q[11318]= 16'he28c;
assign q[11319]= 16'hddce;
assign q[11320]= 16'hd9db;
assign q[11321]= 16'hd6c5;
assign q[11322]= 16'hd496;
assign q[11323]= 16'hd351;
assign q[11324]= 16'hd2ee;
assign q[11325]= 16'hd362;
assign q[11326]= 16'hd498;
assign q[11327]= 16'hd675;
assign q[11328]= 16'hd8dc;
assign q[11329]= 16'hdbab;
assign q[11330]= 16'hdebd;
assign q[11331]= 16'he1ef;
assign q[11332]= 16'he51b;
assign q[11333]= 16'he820;
assign q[11334]= 16'headf;
assign q[11335]= 16'hed3d;
assign q[11336]= 16'hef24;
assign q[11337]= 16'hf084;
assign q[11338]= 16'hf151;
assign q[11339]= 16'hf187;
assign q[11340]= 16'hf127;
assign q[11341]= 16'hf037;
assign q[11342]= 16'heec2;
assign q[11343]= 16'hecd8;
assign q[11344]= 16'hea8c;
assign q[11345]= 16'he7f3;
assign q[11346]= 16'he524;
assign q[11347]= 16'he236;
assign q[11348]= 16'hdf42;
assign q[11349]= 16'hdc5c;
assign q[11350]= 16'hd998;
assign q[11351]= 16'hd708;
assign q[11352]= 16'hd4bb;
assign q[11353]= 16'hd2bb;
assign q[11354]= 16'hd10f;
assign q[11355]= 16'hcfbc;
assign q[11356]= 16'hcec3;
assign q[11357]= 16'hce20;
assign q[11358]= 16'hcdd0;
assign q[11359]= 16'hcdc9;
assign q[11360]= 16'hce04;
assign q[11361]= 16'hce76;
assign q[11362]= 16'hcf14;
assign q[11363]= 16'hcfd3;
assign q[11364]= 16'hd0a8;
assign q[11365]= 16'hd18a;
assign q[11366]= 16'hd26e;
assign q[11367]= 16'hd34e;
assign q[11368]= 16'hd423;
assign q[11369]= 16'hd4e6;
assign q[11370]= 16'hd595;
assign q[11371]= 16'hd62c;
assign q[11372]= 16'hd6a8;
assign q[11373]= 16'hd70a;
assign q[11374]= 16'hd74f;
assign q[11375]= 16'hd778;
assign q[11376]= 16'hd784;
assign q[11377]= 16'hd773;
assign q[11378]= 16'hd746;
assign q[11379]= 16'hd6fd;
assign q[11380]= 16'hd697;
assign q[11381]= 16'hd615;
assign q[11382]= 16'hd577;
assign q[11383]= 16'hd4c0;
assign q[11384]= 16'hd3f1;
assign q[11385]= 16'hd30e;
assign q[11386]= 16'hd21b;
assign q[11387]= 16'hd11f;
assign q[11388]= 16'hd021;
assign q[11389]= 16'hcf2b;
assign q[11390]= 16'hce49;
assign q[11391]= 16'hcd86;
assign q[11392]= 16'hccf1;
assign q[11393]= 16'hcc99;
assign q[11394]= 16'hcc8d;
assign q[11395]= 16'hccdb;
assign q[11396]= 16'hcd94;
assign q[11397]= 16'hcec3;
assign q[11398]= 16'hd074;
assign q[11399]= 16'hd2af;
assign q[11400]= 16'hd57a;
assign q[11401]= 16'hd8d8;
assign q[11402]= 16'hdcc4;
assign q[11403]= 16'he13a;
assign q[11404]= 16'he62e;
assign q[11405]= 16'heb92;
assign q[11406]= 16'hf152;
assign q[11407]= 16'hf757;
assign q[11408]= 16'hfd89;
assign q[11409]= 16'h3ca;
assign q[11410]= 16'ha01;
assign q[11411]= 16'h100e;
assign q[11412]= 16'h15d6;
assign q[11413]= 16'h1b3e;
assign q[11414]= 16'h202d;
assign q[11415]= 16'h2491;
assign q[11416]= 16'h2859;
assign q[11417]= 16'h2b7a;
assign q[11418]= 16'h2df0;
assign q[11419]= 16'h2fbb;
assign q[11420]= 16'h30e1;
assign q[11421]= 16'h316f;
assign q[11422]= 16'h3175;
assign q[11423]= 16'h3109;
assign q[11424]= 16'h3043;
assign q[11425]= 16'h2f3e;
assign q[11426]= 16'h2e15;
assign q[11427]= 16'h2ce6;
assign q[11428]= 16'h2bcb;
assign q[11429]= 16'h2adb;
assign q[11430]= 16'h2a2c;
assign q[11431]= 16'h29cd;
assign q[11432]= 16'h29c8;
assign q[11433]= 16'h2a21;
assign q[11434]= 16'h2ad8;
assign q[11435]= 16'h2be3;
assign q[11436]= 16'h2d33;
assign q[11437]= 16'h2eb5;
assign q[11438]= 16'h3050;
assign q[11439]= 16'h31e8;
assign q[11440]= 16'h335c;
assign q[11441]= 16'h348c;
assign q[11442]= 16'h3559;
assign q[11443]= 16'h35a4;
assign q[11444]= 16'h3551;
assign q[11445]= 16'h3449;
assign q[11446]= 16'h327b;
assign q[11447]= 16'h2fdd;
assign q[11448]= 16'h2c6b;
assign q[11449]= 16'h282a;
assign q[11450]= 16'h2327;
assign q[11451]= 16'h1d76;
assign q[11452]= 16'h1733;
assign q[11453]= 16'h1080;
assign q[11454]= 16'h986;
assign q[11455]= 16'h26f;
assign q[11456]= 16'hfb6d;
assign q[11457]= 16'hf4ac;
assign q[11458]= 16'hee5d;
assign q[11459]= 16'he8ae;
assign q[11460]= 16'he3c6;
assign q[11461]= 16'hdfca;
assign q[11462]= 16'hdcd6;
assign q[11463]= 16'hdb00;
assign q[11464]= 16'hda56;
assign q[11465]= 16'hdad9;
assign q[11466]= 16'hdc86;
assign q[11467]= 16'hdf4e;
assign q[11468]= 16'he319;
assign q[11469]= 16'he7ca;
assign q[11470]= 16'hed3c;
assign q[11471]= 16'hf344;
assign q[11472]= 16'hf9b4;
assign q[11473]= 16'h5b;
assign q[11474]= 16'h70a;
assign q[11475]= 16'hd90;
assign q[11476]= 16'h13c1;
assign q[11477]= 16'h1974;
assign q[11478]= 16'h1e86;
assign q[11479]= 16'h22d9;
assign q[11480]= 16'h265a;
assign q[11481]= 16'h28f9;
assign q[11482]= 16'h2ab3;
assign q[11483]= 16'h2b89;
assign q[11484]= 16'h2b87;
assign q[11485]= 16'h2abe;
assign q[11486]= 16'h2946;
assign q[11487]= 16'h273b;
assign q[11488]= 16'h24bf;
assign q[11489]= 16'h21f4;
assign q[11490]= 16'h1f00;
assign q[11491]= 16'h1c07;
assign q[11492]= 16'h192c;
assign q[11493]= 16'h168f;
assign q[11494]= 16'h144b;
assign q[11495]= 16'h1279;
assign q[11496]= 16'h112a;
assign q[11497]= 16'h106b;
assign q[11498]= 16'h103f;
assign q[11499]= 16'h10a7;
assign q[11500]= 16'h119c;
assign q[11501]= 16'h1310;
assign q[11502]= 16'h14f2;
assign q[11503]= 16'h172c;
assign q[11504]= 16'h19a4;
assign q[11505]= 16'h1c3e;
assign q[11506]= 16'h1edd;
assign q[11507]= 16'h2164;
assign q[11508]= 16'h23b5;
assign q[11509]= 16'h25b6;
assign q[11510]= 16'h274f;
assign q[11511]= 16'h286a;
assign q[11512]= 16'h28f8;
assign q[11513]= 16'h28eb;
assign q[11514]= 16'h283e;
assign q[11515]= 16'h26ed;
assign q[11516]= 16'h24fc;
assign q[11517]= 16'h2272;
assign q[11518]= 16'h1f5b;
assign q[11519]= 16'h1bc8;
assign q[11520]= 16'h17cd;
assign q[11521]= 16'h137e;
assign q[11522]= 16'hef4;
assign q[11523]= 16'ha49;
assign q[11524]= 16'h596;
assign q[11525]= 16'hf5;
assign q[11526]= 16'hfc7e;
assign q[11527]= 16'hf845;
assign q[11528]= 16'hf461;
assign q[11529]= 16'hf0e2;
assign q[11530]= 16'hedd7;
assign q[11531]= 16'heb4a;
assign q[11532]= 16'he943;
assign q[11533]= 16'he7c5;
assign q[11534]= 16'he6d1;
assign q[11535]= 16'he665;
assign q[11536]= 16'he67c;
assign q[11537]= 16'he70c;
assign q[11538]= 16'he80d;
assign q[11539]= 16'he974;
assign q[11540]= 16'heb34;
assign q[11541]= 16'hed41;
assign q[11542]= 16'hef8e;
assign q[11543]= 16'hf210;
assign q[11544]= 16'hf4bc;
assign q[11545]= 16'hf787;
assign q[11546]= 16'hfa68;
assign q[11547]= 16'hfd5b;
assign q[11548]= 16'h57;
assign q[11549]= 16'h35c;
assign q[11550]= 16'h666;
assign q[11551]= 16'h975;
assign q[11552]= 16'hc88;
assign q[11553]= 16'hf9f;
assign q[11554]= 16'h12bc;
assign q[11555]= 16'h15df;
assign q[11556]= 16'h1907;
assign q[11557]= 16'h1c33;
assign q[11558]= 16'h1f61;
assign q[11559]= 16'h228c;
assign q[11560]= 16'h25ae;
assign q[11561]= 16'h28bf;
assign q[11562]= 16'h2bb4;
assign q[11563]= 16'h2e82;
assign q[11564]= 16'h311b;
assign q[11565]= 16'h3370;
assign q[11566]= 16'h3573;
assign q[11567]= 16'h3712;
assign q[11568]= 16'h3840;
assign q[11569]= 16'h38ed;
assign q[11570]= 16'h390f;
assign q[11571]= 16'h3899;
assign q[11572]= 16'h3787;
assign q[11573]= 16'h35d4;
assign q[11574]= 16'h3380;
assign q[11575]= 16'h3092;
assign q[11576]= 16'h2d13;
assign q[11577]= 16'h2911;
assign q[11578]= 16'h249f;
assign q[11579]= 16'h1fd3;
assign q[11580]= 16'h1ac9;
assign q[11581]= 16'h159e;
assign q[11582]= 16'h1071;
assign q[11583]= 16'hb63;
assign q[11584]= 16'h695;
assign q[11585]= 16'h228;
assign q[11586]= 16'hfe3a;
assign q[11587]= 16'hfae5;
assign q[11588]= 16'hf842;
assign q[11589]= 16'hf662;
assign q[11590]= 16'hf553;
assign q[11591]= 16'hf51b;
assign q[11592]= 16'hf5bb;
assign q[11593]= 16'hf72b;
assign q[11594]= 16'hf95f;
assign q[11595]= 16'hfc43;
assign q[11596]= 16'hffbe;
assign q[11597]= 16'h3b0;
assign q[11598]= 16'h7f9;
assign q[11599]= 16'hc73;
assign q[11600]= 16'h10f6;
assign q[11601]= 16'h155b;
assign q[11602]= 16'h197a;
assign q[11603]= 16'h1d2e;
assign q[11604]= 16'h2054;
assign q[11605]= 16'h22d0;
assign q[11606]= 16'h2487;
assign q[11607]= 16'h2568;
assign q[11608]= 16'h2565;
assign q[11609]= 16'h247a;
assign q[11610]= 16'h22a8;
assign q[11611]= 16'h1ff6;
assign q[11612]= 16'h1c73;
assign q[11613]= 16'h1834;
assign q[11614]= 16'h1351;
assign q[11615]= 16'hde8;
assign q[11616]= 16'h819;
assign q[11617]= 16'h209;
assign q[11618]= 16'hfbda;
assign q[11619]= 16'hf5b0;
assign q[11620]= 16'hefad;
assign q[11621]= 16'he9f3;
assign q[11622]= 16'he4a0;
assign q[11623]= 16'hdfcd;
assign q[11624]= 16'hdb91;
assign q[11625]= 16'hd7fd;
assign q[11626]= 16'hd51f;
assign q[11627]= 16'hd2ff;
assign q[11628]= 16'hd1a0;
assign q[11629]= 16'hd101;
assign q[11630]= 16'hd11e;
assign q[11631]= 16'hd1ee;
assign q[11632]= 16'hd365;
assign q[11633]= 16'hd576;
assign q[11634]= 16'hd80f;
assign q[11635]= 16'hdb1f;
assign q[11636]= 16'hde92;
assign q[11637]= 16'he255;
assign q[11638]= 16'he653;
assign q[11639]= 16'hea79;
assign q[11640]= 16'heeb4;
assign q[11641]= 16'hf2ef;
assign q[11642]= 16'hf719;
assign q[11643]= 16'hfb20;
assign q[11644]= 16'hfef5;
assign q[11645]= 16'h285;
assign q[11646]= 16'h5c6;
assign q[11647]= 16'h8a8;
assign q[11648]= 16'hb22;
assign q[11649]= 16'hd28;
assign q[11650]= 16'heb4;
assign q[11651]= 16'hfbe;
assign q[11652]= 16'h1044;
assign q[11653]= 16'h1043;
assign q[11654]= 16'hfbf;
assign q[11655]= 16'hebc;
assign q[11656]= 16'hd40;
assign q[11657]= 16'hb59;
assign q[11658]= 16'h914;
assign q[11659]= 16'h682;
assign q[11660]= 16'h3b7;
assign q[11661]= 16'hcc;
assign q[11662]= 16'hfdd9;
assign q[11663]= 16'hfaf7;
assign q[11664]= 16'hf842;
assign q[11665]= 16'hf5d5;
assign q[11666]= 16'hf3ca;
assign q[11667]= 16'hf23a;
assign q[11668]= 16'hf138;
assign q[11669]= 16'hf0d7;
assign q[11670]= 16'hf122;
assign q[11671]= 16'hf223;
assign q[11672]= 16'hf3d9;
assign q[11673]= 16'hf641;
assign q[11674]= 16'hf94f;
assign q[11675]= 16'hfcf3;
assign q[11676]= 16'h112;
assign q[11677]= 16'h593;
assign q[11678]= 16'ha53;
assign q[11679]= 16'hf2b;
assign q[11680]= 16'h13f6;
assign q[11681]= 16'h1889;
assign q[11682]= 16'h1cbb;
assign q[11683]= 16'h2066;
assign q[11684]= 16'h2365;
assign q[11685]= 16'h2598;
assign q[11686]= 16'h26e7;
assign q[11687]= 16'h273d;
assign q[11688]= 16'h2690;
assign q[11689]= 16'h24dd;
assign q[11690]= 16'h222a;
assign q[11691]= 16'h1e84;
assign q[11692]= 16'h1a03;
assign q[11693]= 16'h14c5;
assign q[11694]= 16'hef0;
assign q[11695]= 16'h8ad;
assign q[11696]= 16'h22c;
assign q[11697]= 16'hfb9f;
assign q[11698]= 16'hf538;
assign q[11699]= 16'hef2a;
assign q[11700]= 16'he9a4;
assign q[11701]= 16'he4d1;
assign q[11702]= 16'he0da;
assign q[11703]= 16'hdddc;
assign q[11704]= 16'hdbf1;
assign q[11705]= 16'hdb28;
assign q[11706]= 16'hdb88;
assign q[11707]= 16'hdd0d;
assign q[11708]= 16'hdfae;
assign q[11709]= 16'he357;
assign q[11710]= 16'he7ec;
assign q[11711]= 16'hed4c;
assign q[11712]= 16'hf350;
assign q[11713]= 16'hf9cd;
assign q[11714]= 16'h95;
assign q[11715]= 16'h77a;
assign q[11716]= 16'he4e;
assign q[11717]= 16'h14e5;
assign q[11718]= 16'h1b15;
assign q[11719]= 16'h20bb;
assign q[11720]= 16'h25b5;
assign q[11721]= 16'h29ec;
assign q[11722]= 16'h2d4b;
assign q[11723]= 16'h2fc6;
assign q[11724]= 16'h3157;
assign q[11725]= 16'h31ff;
assign q[11726]= 16'h31c4;
assign q[11727]= 16'h30b0;
assign q[11728]= 16'h2ed5;
assign q[11729]= 16'h2c45;
assign q[11730]= 16'h2917;
assign q[11731]= 16'h2562;
assign q[11732]= 16'h2141;
assign q[11733]= 16'h1ccc;
assign q[11734]= 16'h181a;
assign q[11735]= 16'h1344;
assign q[11736]= 16'he5d;
assign q[11737]= 16'h979;
assign q[11738]= 16'h4a8;
assign q[11739]= 16'hfff9;
assign q[11740]= 16'hfb74;
assign q[11741]= 16'hf723;
assign q[11742]= 16'hf30e;
assign q[11743]= 16'hef37;
assign q[11744]= 16'heba3;
assign q[11745]= 16'he852;
assign q[11746]= 16'he544;
assign q[11747]= 16'he27a;
assign q[11748]= 16'hdff2;
assign q[11749]= 16'hddab;
assign q[11750]= 16'hdba3;
assign q[11751]= 16'hd9da;
assign q[11752]= 16'hd84d;
assign q[11753]= 16'hd6f9;
assign q[11754]= 16'hd5de;
assign q[11755]= 16'hd4f8;
assign q[11756]= 16'hd445;
assign q[11757]= 16'hd3bf;
assign q[11758]= 16'hd364;
assign q[11759]= 16'hd32d;
assign q[11760]= 16'hd315;
assign q[11761]= 16'hd316;
assign q[11762]= 16'hd327;
assign q[11763]= 16'hd343;
assign q[11764]= 16'hd362;
assign q[11765]= 16'hd37c;
assign q[11766]= 16'hd38b;
assign q[11767]= 16'hd389;
assign q[11768]= 16'hd372;
assign q[11769]= 16'hd344;
assign q[11770]= 16'hd2fd;
assign q[11771]= 16'hd29e;
assign q[11772]= 16'hd22c;
assign q[11773]= 16'hd1ab;
assign q[11774]= 16'hd124;
assign q[11775]= 16'hd0a0;
assign q[11776]= 16'hd02c;
assign q[11777]= 16'hcfd3;
assign q[11778]= 16'hcfa5;
assign q[11779]= 16'hcfae;
assign q[11780]= 16'hcffc;
assign q[11781]= 16'hd09c;
assign q[11782]= 16'hd19a;
assign q[11783]= 16'hd2fc;
assign q[11784]= 16'hd4cb;
assign q[11785]= 16'hd707;
assign q[11786]= 16'hd9b0;
assign q[11787]= 16'hdcc2;
assign q[11788]= 16'he033;
assign q[11789]= 16'he3f7;
assign q[11790]= 16'he7fd;
assign q[11791]= 16'hec34;
assign q[11792]= 16'hf083;
assign q[11793]= 16'hf4d5;
assign q[11794]= 16'hf90f;
assign q[11795]= 16'hfd18;
assign q[11796]= 16'hd7;
assign q[11797]= 16'h438;
assign q[11798]= 16'h723;
assign q[11799]= 16'h988;
assign q[11800]= 16'hb59;
assign q[11801]= 16'hc8e;
assign q[11802]= 16'hd21;
assign q[11803]= 16'hd14;
assign q[11804]= 16'hc6d;
assign q[11805]= 16'hb37;
assign q[11806]= 16'h981;
assign q[11807]= 16'h760;
assign q[11808]= 16'h4e9;
assign q[11809]= 16'h236;
assign q[11810]= 16'hff63;
assign q[11811]= 16'hfc89;
assign q[11812]= 16'hf9c3;
assign q[11813]= 16'hf729;
assign q[11814]= 16'hf4d3;
assign q[11815]= 16'hf2d1;
assign q[11816]= 16'hf132;
assign q[11817]= 16'hefff;
assign q[11818]= 16'hef3b;
assign q[11819]= 16'heee6;
assign q[11820]= 16'heef6;
assign q[11821]= 16'hef62;
assign q[11822]= 16'hf017;
assign q[11823]= 16'hf100;
assign q[11824]= 16'hf208;
assign q[11825]= 16'hf313;
assign q[11826]= 16'hf409;
assign q[11827]= 16'hf4cf;
assign q[11828]= 16'hf54d;
assign q[11829]= 16'hf570;
assign q[11830]= 16'hf525;
assign q[11831]= 16'hf461;
assign q[11832]= 16'hf31d;
assign q[11833]= 16'hf158;
assign q[11834]= 16'hef19;
assign q[11835]= 16'hec6d;
assign q[11836]= 16'he965;
assign q[11837]= 16'he61b;
assign q[11838]= 16'he2ab;
assign q[11839]= 16'hdf37;
assign q[11840]= 16'hdbe2;
assign q[11841]= 16'hd8d1;
assign q[11842]= 16'hd629;
assign q[11843]= 16'hd40e;
assign q[11844]= 16'hd29f;
assign q[11845]= 16'hd1f8;
assign q[11846]= 16'hd22f;
assign q[11847]= 16'hd353;
assign q[11848]= 16'hd56c;
assign q[11849]= 16'hd877;
assign q[11850]= 16'hdc6d;
assign q[11851]= 16'he13b;
assign q[11852]= 16'he6c8;
assign q[11853]= 16'hecf2;
assign q[11854]= 16'hf391;
assign q[11855]= 16'hfa7a;
assign q[11856]= 16'h17b;
assign q[11857]= 16'h865;
assign q[11858]= 16'hf03;
assign q[11859]= 16'h1527;
assign q[11860]= 16'h1aa2;
assign q[11861]= 16'h1f4e;
assign q[11862]= 16'h230a;
assign q[11863]= 16'h25bb;
assign q[11864]= 16'h2753;
assign q[11865]= 16'h27ca;
assign q[11866]= 16'h2725;
assign q[11867]= 16'h2571;
assign q[11868]= 16'h22c4;
assign q[11869]= 16'h1f3e;
assign q[11870]= 16'h1b07;
assign q[11871]= 16'h164b;
assign q[11872]= 16'h113e;
assign q[11873]= 16'hc12;
assign q[11874]= 16'h6fe;
assign q[11875]= 16'h235;
assign q[11876]= 16'hfde9;
assign q[11877]= 16'hfa44;
assign q[11878]= 16'hf76a;
assign q[11879]= 16'hf579;
assign q[11880]= 16'hf484;
assign q[11881]= 16'hf495;
assign q[11882]= 16'hf5aa;
assign q[11883]= 16'hf7b9;
assign q[11884]= 16'hfaad;
assign q[11885]= 16'hfe68;
assign q[11886]= 16'h2c4;
assign q[11887]= 16'h797;
assign q[11888]= 16'hcb0;
assign q[11889]= 16'h11dc;
assign q[11890]= 16'h16e8;
assign q[11891]= 16'h1ba2;
assign q[11892]= 16'h1fdb;
assign q[11893]= 16'h2369;
assign q[11894]= 16'h262a;
assign q[11895]= 16'h2804;
assign q[11896]= 16'h28e4;
assign q[11897]= 16'h28c3;
assign q[11898]= 16'h27a4;
assign q[11899]= 16'h2592;
assign q[11900]= 16'h22a3;
assign q[11901]= 16'h1ef4;
assign q[11902]= 16'h1aab;
assign q[11903]= 16'h15f2;
assign q[11904]= 16'h10f9;
assign q[11905]= 16'hbf0;
assign q[11906]= 16'h709;
assign q[11907]= 16'h273;
assign q[11908]= 16'hfe5b;
assign q[11909]= 16'hfae6;
assign q[11910]= 16'hf836;
assign q[11911]= 16'hf664;
assign q[11912]= 16'hf57f;
assign q[11913]= 16'hf58e;
assign q[11914]= 16'hf68f;
assign q[11915]= 16'hf876;
assign q[11916]= 16'hfb30;
assign q[11917]= 16'hfe9f;
assign q[11918]= 16'h2a1;
assign q[11919]= 16'h70f;
assign q[11920]= 16'hbbd;
assign q[11921]= 16'h107d;
assign q[11922]= 16'h1520;
assign q[11923]= 16'h197a;
assign q[11924]= 16'h1d60;
assign q[11925]= 16'h20ab;
assign q[11926]= 16'h233b;
assign q[11927]= 16'h24f4;
assign q[11928]= 16'h25c4;
assign q[11929]= 16'h259e;
assign q[11930]= 16'h247d;
assign q[11931]= 16'h2266;
assign q[11932]= 16'h1f62;
assign q[11933]= 16'h1b84;
assign q[11934]= 16'h16e2;
assign q[11935]= 16'h1198;
assign q[11936]= 16'hbc9;
assign q[11937]= 16'h596;
assign q[11938]= 16'hff26;
assign q[11939]= 16'hf89c;
assign q[11940]= 16'hf220;
assign q[11941]= 16'hebd5;
assign q[11942]= 16'he5dd;
assign q[11943]= 16'he056;
assign q[11944]= 16'hdb5d;
assign q[11945]= 16'hd707;
assign q[11946]= 16'hd369;
assign q[11947]= 16'hd091;
assign q[11948]= 16'hce89;
assign q[11949]= 16'hcd57;
assign q[11950]= 16'hccfd;
assign q[11951]= 16'hcd7a;
assign q[11952]= 16'hcec6;
assign q[11953]= 16'hd0db;
assign q[11954]= 16'hd3ab;
assign q[11955]= 16'hd728;
assign q[11956]= 16'hdb42;
assign q[11957]= 16'hdfe6;
assign q[11958]= 16'he500;
assign q[11959]= 16'hea78;
assign q[11960]= 16'hf039;
assign q[11961]= 16'hf629;
assign q[11962]= 16'hfc2f;
assign q[11963]= 16'h231;
assign q[11964]= 16'h816;
assign q[11965]= 16'hdc2;
assign q[11966]= 16'h131d;
assign q[11967]= 16'h180d;
assign q[11968]= 16'h1c7a;
assign q[11969]= 16'h204e;
assign q[11970]= 16'h2375;
assign q[11971]= 16'h25de;
assign q[11972]= 16'h277a;
assign q[11973]= 16'h283f;
assign q[11974]= 16'h2828;
assign q[11975]= 16'h2732;
assign q[11976]= 16'h2561;
assign q[11977]= 16'h22bd;
assign q[11978]= 16'h1f54;
assign q[11979]= 16'h1b37;
assign q[11980]= 16'h167e;
assign q[11981]= 16'h1145;
assign q[11982]= 16'hbaa;
assign q[11983]= 16'h5d0;
assign q[11984]= 16'hffdc;
assign q[11985]= 16'hf9f3;
assign q[11986]= 16'hf43b;
assign q[11987]= 16'heeda;
assign q[11988]= 16'he9f5;
assign q[11989]= 16'he5ac;
assign q[11990]= 16'he21e;
assign q[11991]= 16'hdf64;
assign q[11992]= 16'hdd91;
assign q[11993]= 16'hdcb6;
assign q[11994]= 16'hdcd8;
assign q[11995]= 16'hddfc;
assign q[11996]= 16'he01b;
assign q[11997]= 16'he32c;
assign q[11998]= 16'he71d;
assign q[11999]= 16'hebd9;
assign q[12000]= 16'hf144;
assign q[12001]= 16'hf741;
assign q[12002]= 16'hfdad;
assign q[12003]= 16'h464;
assign q[12004]= 16'hb43;
assign q[12005]= 16'h1225;
assign q[12006]= 16'h18e4;
assign q[12007]= 16'h1f60;
assign q[12008]= 16'h2578;
assign q[12009]= 16'h2b10;
assign q[12010]= 16'h300f;
assign q[12011]= 16'h3462;
assign q[12012]= 16'h37f8;
assign q[12013]= 16'h3ac6;
assign q[12014]= 16'h3cc7;
assign q[12015]= 16'h3df8;
assign q[12016]= 16'h3e5b;
assign q[12017]= 16'h3df8;
assign q[12018]= 16'h3cd9;
assign q[12019]= 16'h3b0a;
assign q[12020]= 16'h389c;
assign q[12021]= 16'h35a1;
assign q[12022]= 16'h322b;
assign q[12023]= 16'h2e51;
assign q[12024]= 16'h2a28;
assign q[12025]= 16'h25c5;
assign q[12026]= 16'h213d;
assign q[12027]= 16'h1ca6;
assign q[12028]= 16'h1814;
assign q[12029]= 16'h139a;
assign q[12030]= 16'hf4b;
assign q[12031]= 16'hb37;
assign q[12032]= 16'h76e;
assign q[12033]= 16'h3fd;
assign q[12034]= 16'hf0;
assign q[12035]= 16'hfe54;
assign q[12036]= 16'hfc2f;
assign q[12037]= 16'hfa88;
assign q[12038]= 16'hf965;
assign q[12039]= 16'hf8c8;
assign q[12040]= 16'hf8b3;
assign q[12041]= 16'hf925;
assign q[12042]= 16'hfa1b;
assign q[12043]= 16'hfb8f;
assign q[12044]= 16'hfd7b;
assign q[12045]= 16'hffd4;
assign q[12046]= 16'h290;
assign q[12047]= 16'h5a2;
assign q[12048]= 16'h8fc;
assign q[12049]= 16'hc8d;
assign q[12050]= 16'h1043;
assign q[12051]= 16'h140c;
assign q[12052]= 16'h17d6;
assign q[12053]= 16'h1b8d;
assign q[12054]= 16'h1f1c;
assign q[12055]= 16'h2272;
assign q[12056]= 16'h257c;
assign q[12057]= 16'h2829;
assign q[12058]= 16'h2a68;
assign q[12059]= 16'h2c2d;
assign q[12060]= 16'h2d6b;
assign q[12061]= 16'h2e17;
assign q[12062]= 16'h2e2c;
assign q[12063]= 16'h2da5;
assign q[12064]= 16'h2c7f;
assign q[12065]= 16'h2abd;
assign q[12066]= 16'h2861;
assign q[12067]= 16'h2573;
assign q[12068]= 16'h21fb;
assign q[12069]= 16'h1e07;
assign q[12070]= 16'h19a4;
assign q[12071]= 16'h14e2;
assign q[12072]= 16'hfd5;
assign q[12073]= 16'ha90;
assign q[12074]= 16'h528;
assign q[12075]= 16'hffb6;
assign q[12076]= 16'hfa4f;
assign q[12077]= 16'hf509;
assign q[12078]= 16'heffe;
assign q[12079]= 16'heb44;
assign q[12080]= 16'he6f0;
assign q[12081]= 16'he316;
assign q[12082]= 16'hdfcb;
assign q[12083]= 16'hdd1e;
assign q[12084]= 16'hdb1d;
assign q[12085]= 16'hd9d5;
assign q[12086]= 16'hd94c;
assign q[12087]= 16'hd987;
assign q[12088]= 16'hda89;
assign q[12089]= 16'hdc4e;
assign q[12090]= 16'hded0;
assign q[12091]= 16'he204;
assign q[12092]= 16'he5de;
assign q[12093]= 16'hea4b;
assign q[12094]= 16'hef39;
assign q[12095]= 16'hf48f;
assign q[12096]= 16'hfa36;
assign q[12097]= 16'h11;
assign q[12098]= 16'h607;
assign q[12099]= 16'hbfc;
assign q[12100]= 16'h11d4;
assign q[12101]= 16'h1775;
assign q[12102]= 16'h1cc6;
assign q[12103]= 16'h21b2;
assign q[12104]= 16'h2626;
assign q[12105]= 16'h2a13;
assign q[12106]= 16'h2d6e;
assign q[12107]= 16'h302f;
assign q[12108]= 16'h3254;
assign q[12109]= 16'h33de;
assign q[12110]= 16'h34d3;
assign q[12111]= 16'h353c;
assign q[12112]= 16'h3525;
assign q[12113]= 16'h349e;
assign q[12114]= 16'h33b7;
assign q[12115]= 16'h3285;
assign q[12116]= 16'h3118;
assign q[12117]= 16'h2f85;
assign q[12118]= 16'h2ddc;
assign q[12119]= 16'h2c2f;
assign q[12120]= 16'h2a89;
assign q[12121]= 16'h28f5;
assign q[12122]= 16'h277b;
assign q[12123]= 16'h261e;
assign q[12124]= 16'h24dd;
assign q[12125]= 16'h23b5;
assign q[12126]= 16'h229e;
assign q[12127]= 16'h2190;
assign q[12128]= 16'h207d;
assign q[12129]= 16'h1f58;
assign q[12130]= 16'h1e11;
assign q[12131]= 16'h1c9b;
assign q[12132]= 16'h1ae7;
assign q[12133]= 16'h18e8;
assign q[12134]= 16'h1695;
assign q[12135]= 16'h13e7;
assign q[12136]= 16'h10da;
assign q[12137]= 16'hd6f;
assign q[12138]= 16'h9ab;
assign q[12139]= 16'h596;
assign q[12140]= 16'h13d;
assign q[12141]= 16'hfcb3;
assign q[12142]= 16'hf808;
assign q[12143]= 16'hf355;
assign q[12144]= 16'heeb2;
assign q[12145]= 16'hea38;
assign q[12146]= 16'he600;
assign q[12147]= 16'he221;
assign q[12148]= 16'hdeb3;
assign q[12149]= 16'hdbc7;
assign q[12150]= 16'hd96e;
assign q[12151]= 16'hd7b2;
assign q[12152]= 16'hd699;
assign q[12153]= 16'hd625;
assign q[12154]= 16'hd652;
assign q[12155]= 16'hd715;
assign q[12156]= 16'hd862;
assign q[12157]= 16'hda24;
assign q[12158]= 16'hdc45;
assign q[12159]= 16'hdead;
assign q[12160]= 16'he13f;
assign q[12161]= 16'he3df;
assign q[12162]= 16'he670;
assign q[12163]= 16'he8d8;
assign q[12164]= 16'heafd;
assign q[12165]= 16'hecc8;
assign q[12166]= 16'hee28;
assign q[12167]= 16'hef0e;
assign q[12168]= 16'hef72;
assign q[12169]= 16'hef50;
assign q[12170]= 16'heea9;
assign q[12171]= 16'hed85;
assign q[12172]= 16'hebf0;
assign q[12173]= 16'he9fb;
assign q[12174]= 16'he7ba;
assign q[12175]= 16'he545;
assign q[12176]= 16'he2b7;
assign q[12177]= 16'he02a;
assign q[12178]= 16'hddbb;
assign q[12179]= 16'hdb83;
assign q[12180]= 16'hd99d;
assign q[12181]= 16'hd81f;
assign q[12182]= 16'hd71c;
assign q[12183]= 16'hd6a4;
assign q[12184]= 16'hd6c2;
assign q[12185]= 16'hd77c;
assign q[12186]= 16'hd8d3;
assign q[12187]= 16'hdac3;
assign q[12188]= 16'hdd44;
assign q[12189]= 16'he048;
assign q[12190]= 16'he3c0;
assign q[12191]= 16'he796;
assign q[12192]= 16'hebb4;
assign q[12193]= 16'hf003;
assign q[12194]= 16'hf468;
assign q[12195]= 16'hf8cb;
assign q[12196]= 16'hfd13;
assign q[12197]= 16'h128;
assign q[12198]= 16'h4f8;
assign q[12199]= 16'h870;
assign q[12200]= 16'hb83;
assign q[12201]= 16'he24;
assign q[12202]= 16'h104f;
assign q[12203]= 16'h1200;
assign q[12204]= 16'h1339;
assign q[12205]= 16'h13ff;
assign q[12206]= 16'h145c;
assign q[12207]= 16'h145a;
assign q[12208]= 16'h1408;
assign q[12209]= 16'h1375;
assign q[12210]= 16'h12b4;
assign q[12211]= 16'h11d4;
assign q[12212]= 16'h10e7;
assign q[12213]= 16'hffd;
assign q[12214]= 16'hf25;
assign q[12215]= 16'he6b;
assign q[12216]= 16'hdd9;
assign q[12217]= 16'hd76;
assign q[12218]= 16'hd45;
assign q[12219]= 16'hd47;
assign q[12220]= 16'hd79;
assign q[12221]= 16'hdd5;
assign q[12222]= 16'he53;
assign q[12223]= 16'hee8;
assign q[12224]= 16'hf87;
assign q[12225]= 16'h1022;
assign q[12226]= 16'h10aa;
assign q[12227]= 16'h1110;
assign q[12228]= 16'h1148;
assign q[12229]= 16'h1143;
assign q[12230]= 16'h10f8;
assign q[12231]= 16'h105e;
assign q[12232]= 16'hf72;
assign q[12233]= 16'he30;
assign q[12234]= 16'hc9b;
assign q[12235]= 16'hab9;
assign q[12236]= 16'h892;
assign q[12237]= 16'h634;
assign q[12238]= 16'h3ad;
assign q[12239]= 16'h110;
assign q[12240]= 16'hfe71;
assign q[12241]= 16'hfbe2;
assign q[12242]= 16'hf97a;
assign q[12243]= 16'hf74d;
assign q[12244]= 16'hf56f;
assign q[12245]= 16'hf3f0;
assign q[12246]= 16'hf2df;
assign q[12247]= 16'hf246;
assign q[12248]= 16'hf22d;
assign q[12249]= 16'hf294;
assign q[12250]= 16'hf37a;
assign q[12251]= 16'hf4d8;
assign q[12252]= 16'hf6a1;
assign q[12253]= 16'hf8c6;
assign q[12254]= 16'hfb32;
assign q[12255]= 16'hfdd0;
assign q[12256]= 16'h85;
assign q[12257]= 16'h339;
assign q[12258]= 16'h5d0;
assign q[12259]= 16'h831;
assign q[12260]= 16'ha43;
assign q[12261]= 16'hbf1;
assign q[12262]= 16'hd29;
assign q[12263]= 16'hddf;
assign q[12264]= 16'he08;
assign q[12265]= 16'hda4;
assign q[12266]= 16'hcb4;
assign q[12267]= 16'hb41;
assign q[12268]= 16'h959;
assign q[12269]= 16'h70e;
assign q[12270]= 16'h478;
assign q[12271]= 16'h1b0;
assign q[12272]= 16'hfed4;
assign q[12273]= 16'hfc01;
assign q[12274]= 16'hf954;
assign q[12275]= 16'hf6eb;
assign q[12276]= 16'hf4df;
assign q[12277]= 16'hf348;
assign q[12278]= 16'hf238;
assign q[12279]= 16'hf1bb;
assign q[12280]= 16'hf1d8;
assign q[12281]= 16'hf28f;
assign q[12282]= 16'hf3da;
assign q[12283]= 16'hf5ad;
assign q[12284]= 16'hf7f5;
assign q[12285]= 16'hfa9a;
assign q[12286]= 16'hfd80;
assign q[12287]= 16'h85;
