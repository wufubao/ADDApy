assign i[0]= 16'hdc0e;
assign i[1]= 16'hda83;
assign i[2]= 16'hd934;
assign i[3]= 16'hd81e;
assign i[4]= 16'hd738;
assign i[5]= 16'hd67e;
assign i[6]= 16'hd5ea;
assign i[7]= 16'hd574;
assign i[8]= 16'hd51a;
assign i[9]= 16'hd4d4;
assign i[10]= 16'hd49f;
assign i[11]= 16'hd478;
assign i[12]= 16'hd45a;
assign i[13]= 16'hd444;
assign i[14]= 16'hd432;
assign i[15]= 16'hd421;
assign i[16]= 16'hd410;
assign i[17]= 16'hd3fd;
assign i[18]= 16'hd3e5;
assign i[19]= 16'hd3c7;
assign i[20]= 16'hd3a0;
assign i[21]= 16'hd36f;
assign i[22]= 16'hd333;
assign i[23]= 16'hd2ea;
assign i[24]= 16'hd296;
assign i[25]= 16'hd235;
assign i[26]= 16'hd1ca;
assign i[27]= 16'hd158;
assign i[28]= 16'hd0e1;
assign i[29]= 16'hd06b;
assign i[30]= 16'hcffb;
assign i[31]= 16'hcf98;
assign i[32]= 16'hcf49;
assign i[33]= 16'hcf16;
assign i[34]= 16'hcf06;
assign i[35]= 16'hcf22;
assign i[36]= 16'hcf71;
assign i[37]= 16'hcff8;
assign i[38]= 16'hd0be;
assign i[39]= 16'hd1c5;
assign i[40]= 16'hd30e;
assign i[41]= 16'hd498;
assign i[42]= 16'hd660;
assign i[43]= 16'hd860;
assign i[44]= 16'hda8e;
assign i[45]= 16'hdce1;
assign i[46]= 16'hdf4a;
assign i[47]= 16'he1ba;
assign i[48]= 16'he423;
assign i[49]= 16'he671;
assign i[50]= 16'he895;
assign i[51]= 16'hea7e;
assign i[52]= 16'hec1b;
assign i[53]= 16'hed60;
assign i[54]= 16'hee41;
assign i[55]= 16'heeb5;
assign i[56]= 16'heeb8;
assign i[57]= 16'hee48;
assign i[58]= 16'hed68;
assign i[59]= 16'hec1f;
assign i[60]= 16'hea78;
assign i[61]= 16'he881;
assign i[62]= 16'he64b;
assign i[63]= 16'he3eb;
assign i[64]= 16'he178;
assign i[65]= 16'hdf09;
assign i[66]= 16'hdcb7;
assign i[67]= 16'hda9a;
assign i[68]= 16'hd8c9;
assign i[69]= 16'hd75a;
assign i[70]= 16'hd65f;
assign i[71]= 16'hd5e8;
assign i[72]= 16'hd600;
assign i[73]= 16'hd6ae;
assign i[74]= 16'hd7f5;
assign i[75]= 16'hd9d3;
assign i[76]= 16'hdc42;
assign i[77]= 16'hdf36;
assign i[78]= 16'he2a2;
assign i[79]= 16'he673;
assign i[80]= 16'hea94;
assign i[81]= 16'heeee;
assign i[82]= 16'hf369;
assign i[83]= 16'hf7ed;
assign i[84]= 16'hfc60;
assign i[85]= 16'hac;
assign i[86]= 16'h4bb;
assign i[87]= 16'h87b;
assign i[88]= 16'hbdc;
assign i[89]= 16'hed0;
assign i[90]= 16'h114f;
assign i[91]= 16'h1353;
assign i[92]= 16'h14db;
assign i[93]= 16'h15ea;
assign i[94]= 16'h1684;
assign i[95]= 16'h16b1;
assign i[96]= 16'h167c;
assign i[97]= 16'h15f2;
assign i[98]= 16'h151e;
assign i[99]= 16'h1411;
assign i[100]= 16'h12d7;
assign i[101]= 16'h117d;
assign i[102]= 16'h1010;
assign i[103]= 16'he99;
assign i[104]= 16'hd22;
assign i[105]= 16'hbb1;
assign i[106]= 16'ha49;
assign i[107]= 16'h8ec;
assign i[108]= 16'h799;
assign i[109]= 16'h64d;
assign i[110]= 16'h504;
assign i[111]= 16'h3b7;
assign i[112]= 16'h25f;
assign i[113]= 16'hf6;
assign i[114]= 16'hff75;
assign i[115]= 16'hfdd2;
assign i[116]= 16'hfc0a;
assign i[117]= 16'hfa17;
assign i[118]= 16'hf7f7;
assign i[119]= 16'hf5aa;
assign i[120]= 16'hf332;
assign i[121]= 16'hf092;
assign i[122]= 16'hedd2;
assign i[123]= 16'heaf9;
assign i[124]= 16'he815;
assign i[125]= 16'he530;
assign i[126]= 16'he25a;
assign i[127]= 16'hdfa2;
assign i[128]= 16'hdd17;
assign i[129]= 16'hdacb;
assign i[130]= 16'hd8ca;
assign i[131]= 16'hd726;
assign i[132]= 16'hd5e9;
assign i[133]= 16'hd51e;
assign i[134]= 16'hd4cf;
assign i[135]= 16'hd501;
assign i[136]= 16'hd5b8;
assign i[137]= 16'hd6f2;
assign i[138]= 16'hd8ae;
assign i[139]= 16'hdae5;
assign i[140]= 16'hdd90;
assign i[141]= 16'he0a2;
assign i[142]= 16'he410;
assign i[143]= 16'he7ca;
assign i[144]= 16'hebc1;
assign i[145]= 16'hefe3;
assign i[146]= 16'hf420;
assign i[147]= 16'hf868;
assign i[148]= 16'hfcaa;
assign i[149]= 16'hd7;
assign i[150]= 16'h4e3;
assign i[151]= 16'h8c3;
assign i[152]= 16'hc6e;
assign i[153]= 16'hfdc;
assign i[154]= 16'h1309;
assign i[155]= 16'h15f3;
assign i[156]= 16'h189a;
assign i[157]= 16'h1b00;
assign i[158]= 16'h1d2a;
assign i[159]= 16'h1f1c;
assign i[160]= 16'h20dc;
assign i[161]= 16'h2272;
assign i[162]= 16'h23e5;
assign i[163]= 16'h253c;
assign i[164]= 16'h267d;
assign i[165]= 16'h27af;
assign i[166]= 16'h28d5;
assign i[167]= 16'h29f3;
assign i[168]= 16'h2b0b;
assign i[169]= 16'h2c1c;
assign i[170]= 16'h2d24;
assign i[171]= 16'h2e22;
assign i[172]= 16'h2f0f;
assign i[173]= 16'h2fe6;
assign i[174]= 16'h30a1;
assign i[175]= 16'h3137;
assign i[176]= 16'h31a1;
assign i[177]= 16'h31d7;
assign i[178]= 16'h31d2;
assign i[179]= 16'h318a;
assign i[180]= 16'h30fb;
assign i[181]= 16'h301e;
assign i[182]= 16'h2ef2;
assign i[183]= 16'h2d73;
assign i[184]= 16'h2ba2;
assign i[185]= 16'h2981;
assign i[186]= 16'h2712;
assign i[187]= 16'h2459;
assign i[188]= 16'h215d;
assign i[189]= 16'h1e25;
assign i[190]= 16'h1ab7;
assign i[191]= 16'h171d;
assign i[192]= 16'h1360;
assign i[193]= 16'hf88;
assign i[194]= 16'hb9f;
assign i[195]= 16'h7ad;
assign i[196]= 16'h3ba;
assign i[197]= 16'hffd1;
assign i[198]= 16'hfbf5;
assign i[199]= 16'hf82e;
assign i[200]= 16'hf483;
assign i[201]= 16'hf0f9;
assign i[202]= 16'hed93;
assign i[203]= 16'hea57;
assign i[204]= 16'he748;
assign i[205]= 16'he46a;
assign i[206]= 16'he1be;
assign i[207]= 16'hdf48;
assign i[208]= 16'hdd0a;
assign i[209]= 16'hdb05;
assign i[210]= 16'hd93c;
assign i[211]= 16'hd7af;
assign i[212]= 16'hd65f;
assign i[213]= 16'hd54b;
assign i[214]= 16'hd474;
assign i[215]= 16'hd3d7;
assign i[216]= 16'hd371;
assign i[217]= 16'hd33e;
assign i[218]= 16'hd33a;
assign i[219]= 16'hd35e;
assign i[220]= 16'hd3a3;
assign i[221]= 16'hd3ff;
assign i[222]= 16'hd46b;
assign i[223]= 16'hd4dc;
assign i[224]= 16'hd547;
assign i[225]= 16'hd5a4;
assign i[226]= 16'hd5e6;
assign i[227]= 16'hd607;
assign i[228]= 16'hd5fe;
assign i[229]= 16'hd5c5;
assign i[230]= 16'hd559;
assign i[231]= 16'hd4b8;
assign i[232]= 16'hd3e3;
assign i[233]= 16'hd2e0;
assign i[234]= 16'hd1b6;
assign i[235]= 16'hd06f;
assign i[236]= 16'hcf18;
assign i[237]= 16'hcdc2;
assign i[238]= 16'hcc7e;
assign i[239]= 16'hcb61;
assign i[240]= 16'hca7e;
assign i[241]= 16'hc9eb;
assign i[242]= 16'hc9bc;
assign i[243]= 16'hca03;
assign i[244]= 16'hcad2;
assign i[245]= 16'hcc37;
assign i[246]= 16'hce3b;
assign i[247]= 16'hd0e5;
assign i[248]= 16'hd437;
assign i[249]= 16'hd82d;
assign i[250]= 16'hdcbd;
assign i[251]= 16'he1db;
assign i[252]= 16'he773;
assign i[253]= 16'hed6f;
assign i[254]= 16'hf3b4;
assign i[255]= 16'hfa24;
assign i[256]= 16'h9e;
assign i[257]= 16'h702;
assign i[258]= 16'hd2f;
assign i[259]= 16'h1304;
assign i[260]= 16'h1864;
assign i[261]= 16'h1d33;
assign i[262]= 16'h215a;
assign i[263]= 16'h24c9;
assign i[264]= 16'h2771;
assign i[265]= 16'h294e;
assign i[266]= 16'h2a60;
assign i[267]= 16'h2aab;
assign i[268]= 16'h2a3d;
assign i[269]= 16'h2927;
assign i[270]= 16'h2780;
assign i[271]= 16'h2562;
assign i[272]= 16'h22ed;
assign i[273]= 16'h203f;
assign i[274]= 16'h1d79;
assign i[275]= 16'h1abd;
assign i[276]= 16'h1829;
assign i[277]= 16'h15da;
assign i[278]= 16'h13e9;
assign i[279]= 16'h126a;
assign i[280]= 16'h116d;
assign i[281]= 16'h10fa;
assign i[282]= 16'h1117;
assign i[283]= 16'h11c1;
assign i[284]= 16'h12f0;
assign i[285]= 16'h1495;
assign i[286]= 16'h16a0;
assign i[287]= 16'h18f8;
assign i[288]= 16'h1b86;
assign i[289]= 16'h1e2b;
assign i[290]= 16'h20cd;
assign i[291]= 16'h234c;
assign i[292]= 16'h258d;
assign i[293]= 16'h2776;
assign i[294]= 16'h28ef;
assign i[295]= 16'h29e4;
assign i[296]= 16'h2a46;
assign i[297]= 16'h2a0b;
assign i[298]= 16'h292b;
assign i[299]= 16'h27a8;
assign i[300]= 16'h2585;
assign i[301]= 16'h22cb;
assign i[302]= 16'h1f88;
assign i[303]= 16'h1bcc;
assign i[304]= 16'h17ab;
assign i[305]= 16'h133c;
assign i[306]= 16'he94;
assign i[307]= 16'h9cd;
assign i[308]= 16'h4fe;
assign i[309]= 16'h3b;
assign i[310]= 16'hfb9c;
assign i[311]= 16'hf72f;
assign i[312]= 16'hf304;
assign i[313]= 16'hef27;
assign i[314]= 16'heba0;
assign i[315]= 16'he873;
assign i[316]= 16'he5a2;
assign i[317]= 16'he32a;
assign i[318]= 16'he106;
assign i[319]= 16'hdf30;
assign i[320]= 16'hdd9d;
assign i[321]= 16'hdc44;
assign i[322]= 16'hdb18;
assign i[323]= 16'hda0f;
assign i[324]= 16'hd91e;
assign i[325]= 16'hd83a;
assign i[326]= 16'hd75c;
assign i[327]= 16'hd67c;
assign i[328]= 16'hd597;
assign i[329]= 16'hd4aa;
assign i[330]= 16'hd3b5;
assign i[331]= 16'hd2bd;
assign i[332]= 16'hd1c4;
assign i[333]= 16'hd0d4;
assign i[334]= 16'hcff4;
assign i[335]= 16'hcf2e;
assign i[336]= 16'hce8e;
assign i[337]= 16'hce1e;
assign i[338]= 16'hcdeb;
assign i[339]= 16'hcdff;
assign i[340]= 16'hce63;
assign i[341]= 16'hcf1f;
assign i[342]= 16'hd03a;
assign i[343]= 16'hd1b8;
assign i[344]= 16'hd39b;
assign i[345]= 16'hd5e1;
assign i[346]= 16'hd887;
assign i[347]= 16'hdb87;
assign i[348]= 16'hded8;
assign i[349]= 16'he271;
assign i[350]= 16'he643;
assign i[351]= 16'hea41;
assign i[352]= 16'hee5c;
assign i[353]= 16'hf283;
assign i[354]= 16'hf6a5;
assign i[355]= 16'hfab3;
assign i[356]= 16'hfe9c;
assign i[357]= 16'h252;
assign i[358]= 16'h5c8;
assign i[359]= 16'h8f3;
assign i[360]= 16'hbc9;
assign i[361]= 16'he43;
assign i[362]= 16'h105b;
assign i[363]= 16'h1210;
assign i[364]= 16'h1362;
assign i[365]= 16'h1452;
assign i[366]= 16'h14e5;
assign i[367]= 16'h1520;
assign i[368]= 16'h150b;
assign i[369]= 16'h14ae;
assign i[370]= 16'h1413;
assign i[371]= 16'h1343;
assign i[372]= 16'h1247;
assign i[373]= 16'h1129;
assign i[374]= 16'hff1;
assign i[375]= 16'hea7;
assign i[376]= 16'hd50;
assign i[377]= 16'hbf2;
assign i[378]= 16'ha90;
assign i[379]= 16'h92d;
assign i[380]= 16'h7c7;
assign i[381]= 16'h661;
assign i[382]= 16'h4f6;
assign i[383]= 16'h386;
assign i[384]= 16'h20d;
assign i[385]= 16'h89;
assign i[386]= 16'hfef8;
assign i[387]= 16'hfd55;
assign i[388]= 16'hfba1;
assign i[389]= 16'hf9dc;
assign i[390]= 16'hf808;
assign i[391]= 16'hf627;
assign i[392]= 16'hf43e;
assign i[393]= 16'hf255;
assign i[394]= 16'hf074;
assign i[395]= 16'heea5;
assign i[396]= 16'hecf3;
assign i[397]= 16'heb6a;
assign i[398]= 16'hea18;
assign i[399]= 16'he90a;
assign i[400]= 16'he84d;
assign i[401]= 16'he7ec;
assign i[402]= 16'he7f4;
assign i[403]= 16'he86c;
assign i[404]= 16'he95b;
assign i[405]= 16'heac6;
assign i[406]= 16'hecae;
assign i[407]= 16'hef11;
assign i[408]= 16'hf1e8;
assign i[409]= 16'hf52c;
assign i[410]= 16'hf8d1;
assign i[411]= 16'hfcc6;
assign i[412]= 16'hfa;
assign i[413]= 16'h55a;
assign i[414]= 16'h9ce;
assign i[415]= 16'he3f;
assign i[416]= 16'h1296;
assign i[417]= 16'h16b9;
assign i[418]= 16'h1a91;
assign i[419]= 16'h1e08;
assign i[420]= 16'h210a;
assign i[421]= 16'h2384;
assign i[422]= 16'h256a;
assign i[423]= 16'h26ae;
assign i[424]= 16'h274a;
assign i[425]= 16'h273b;
assign i[426]= 16'h2682;
assign i[427]= 16'h2522;
assign i[428]= 16'h2326;
assign i[429]= 16'h2099;
assign i[430]= 16'h1d8a;
assign i[431]= 16'h1a0d;
assign i[432]= 16'h1636;
assign i[433]= 16'h121c;
assign i[434]= 16'hdd5;
assign i[435]= 16'h979;
assign i[436]= 16'h520;
assign i[437]= 16'he1;
assign i[438]= 16'hfcd1;
assign i[439]= 16'hf901;
assign i[440]= 16'hf582;
assign i[441]= 16'hf264;
assign i[442]= 16'hefaf;
assign i[443]= 16'hed6c;
assign i[444]= 16'heb9e;
assign i[445]= 16'hea47;
assign i[446]= 16'he963;
assign i[447]= 16'he8ee;
assign i[448]= 16'he8de;
assign i[449]= 16'he92b;
assign i[450]= 16'he9c7;
assign i[451]= 16'heaa5;
assign i[452]= 16'hebb6;
assign i[453]= 16'heceb;
assign i[454]= 16'hee35;
assign i[455]= 16'hef86;
assign i[456]= 16'hf0cf;
assign i[457]= 16'hf205;
assign i[458]= 16'hf31c;
assign i[459]= 16'hf40b;
assign i[460]= 16'hf4cb;
assign i[461]= 16'hf557;
assign i[462]= 16'hf5ac;
assign i[463]= 16'hf5c9;
assign i[464]= 16'hf5b1;
assign i[465]= 16'hf565;
assign i[466]= 16'hf4eb;
assign i[467]= 16'hf44a;
assign i[468]= 16'hf387;
assign i[469]= 16'hf2ac;
assign i[470]= 16'hf1c2;
assign i[471]= 16'hf0d2;
assign i[472]= 16'hefe4;
assign i[473]= 16'hef01;
assign i[474]= 16'hee32;
assign i[475]= 16'hed7e;
assign i[476]= 16'hecec;
assign i[477]= 16'hec80;
assign i[478]= 16'hec41;
assign i[479]= 16'hec31;
assign i[480]= 16'hec52;
assign i[481]= 16'heca8;
assign i[482]= 16'hed31;
assign i[483]= 16'hedf0;
assign i[484]= 16'heee2;
assign i[485]= 16'hf009;
assign i[486]= 16'hf162;
assign i[487]= 16'hf2ee;
assign i[488]= 16'hf4ab;
assign i[489]= 16'hf698;
assign i[490]= 16'hf8b6;
assign i[491]= 16'hfb03;
assign i[492]= 16'hfd80;
assign i[493]= 16'h2a;
assign i[494]= 16'h305;
assign i[495]= 16'h60e;
assign i[496]= 16'h943;
assign i[497]= 16'hca2;
assign i[498]= 16'h102a;
assign i[499]= 16'h13d4;
assign i[500]= 16'h179b;
assign i[501]= 16'h1b77;
assign i[502]= 16'h1f60;
assign i[503]= 16'h234b;
assign i[504]= 16'h2729;
assign i[505]= 16'h2aed;
assign i[506]= 16'h2e86;
assign i[507]= 16'h31e4;
assign i[508]= 16'h34f3;
assign i[509]= 16'h37a1;
assign i[510]= 16'h39db;
assign i[511]= 16'h3b8f;
assign i[512]= 16'h3cac;
assign i[513]= 16'h3d24;
assign i[514]= 16'h3ce9;
assign i[515]= 16'h3bf3;
assign i[516]= 16'h3a3b;
assign i[517]= 16'h37c0;
assign i[518]= 16'h3484;
assign i[519]= 16'h308e;
assign i[520]= 16'h2beb;
assign i[521]= 16'h26aa;
assign i[522]= 16'h20e1;
assign i[523]= 16'h1aaa;
assign i[524]= 16'h1420;
assign i[525]= 16'hd64;
assign i[526]= 16'h697;
assign i[527]= 16'hffdf;
assign i[528]= 16'hf95e;
assign i[529]= 16'hf337;
assign i[530]= 16'hed8d;
assign i[531]= 16'he880;
assign i[532]= 16'he42c;
assign i[533]= 16'he0aa;
assign i[534]= 16'hde0c;
assign i[535]= 16'hdc63;
assign i[536]= 16'hdbb5;
assign i[537]= 16'hdc07;
assign i[538]= 16'hdd53;
assign i[539]= 16'hdf92;
assign i[540]= 16'he2b4;
assign i[541]= 16'he6a5;
assign i[542]= 16'heb4d;
assign i[543]= 16'hf08f;
assign i[544]= 16'hf64d;
assign i[545]= 16'hfc66;
assign i[546]= 16'h2b6;
assign i[547]= 16'h91d;
assign i[548]= 16'hf79;
assign i[549]= 16'h15a9;
assign i[550]= 16'h1b92;
assign i[551]= 16'h2118;
assign i[552]= 16'h2626;
assign i[553]= 16'h2aaa;
assign i[554]= 16'h2e95;
assign i[555]= 16'h31df;
assign i[556]= 16'h3484;
assign i[557]= 16'h3683;
assign i[558]= 16'h37e0;
assign i[559]= 16'h38a3;
assign i[560]= 16'h38d8;
assign i[561]= 16'h388c;
assign i[562]= 16'h37d0;
assign i[563]= 16'h36b5;
assign i[564]= 16'h354f;
assign i[565]= 16'h33b0;
assign i[566]= 16'h31ec;
assign i[567]= 16'h3015;
assign i[568]= 16'h2e3e;
assign i[569]= 16'h2c77;
assign i[570]= 16'h2acd;
assign i[571]= 16'h294f;
assign i[572]= 16'h2807;
assign i[573]= 16'h26fd;
assign i[574]= 16'h2639;
assign i[575]= 16'h25bd;
assign i[576]= 16'h258d;
assign i[577]= 16'h25a9;
assign i[578]= 16'h260d;
assign i[579]= 16'h26b8;
assign i[580]= 16'h27a2;
assign i[581]= 16'h28c6;
assign i[582]= 16'h2a19;
assign i[583]= 16'h2b92;
assign i[584]= 16'h2d25;
assign i[585]= 16'h2ec7;
assign i[586]= 16'h3069;
assign i[587]= 16'h31fe;
assign i[588]= 16'h3376;
assign i[589]= 16'h34c4;
assign i[590]= 16'h35d9;
assign i[591]= 16'h36a5;
assign i[592]= 16'h371c;
assign i[593]= 16'h3730;
assign i[594]= 16'h36d6;
assign i[595]= 16'h3604;
assign i[596]= 16'h34b1;
assign i[597]= 16'h32d9;
assign i[598]= 16'h3078;
assign i[599]= 16'h2d8e;
assign i[600]= 16'h2a1d;
assign i[601]= 16'h262c;
assign i[602]= 16'h21c2;
assign i[603]= 16'h1cec;
assign i[604]= 16'h17b9;
assign i[605]= 16'h1239;
assign i[606]= 16'hc81;
assign i[607]= 16'h6a5;
assign i[608]= 16'hbc;
assign i[609]= 16'hfae0;
assign i[610]= 16'hf526;
assign i[611]= 16'hefa6;
assign i[612]= 16'hea77;
assign i[613]= 16'he5ae;
assign i[614]= 16'he15e;
assign i[615]= 16'hdd96;
assign i[616]= 16'hda66;
assign i[617]= 16'hd7d5;
assign i[618]= 16'hd5ea;
assign i[619]= 16'hd4a8;
assign i[620]= 16'hd40d;
assign i[621]= 16'hd415;
assign i[622]= 16'hd4b6;
assign i[623]= 16'hd5e6;
assign i[624]= 16'hd795;
assign i[625]= 16'hd9b2;
assign i[626]= 16'hdc2b;
assign i[627]= 16'hdeec;
assign i[628]= 16'he1df;
assign i[629]= 16'he4f0;
assign i[630]= 16'he809;
assign i[631]= 16'heb16;
assign i[632]= 16'hee04;
assign i[633]= 16'hf0c2;
assign i[634]= 16'hf340;
assign i[635]= 16'hf572;
assign i[636]= 16'hf74c;
assign i[637]= 16'hf8c6;
assign i[638]= 16'hf9d9;
assign i[639]= 16'hfa84;
assign i[640]= 16'hfac4;
assign i[641]= 16'hfa9b;
assign i[642]= 16'hfa0c;
assign i[643]= 16'hf91d;
assign i[644]= 16'hf7d4;
assign i[645]= 16'hf63a;
assign i[646]= 16'hf458;
assign i[647]= 16'hf239;
assign i[648]= 16'hefe9;
assign i[649]= 16'hed73;
assign i[650]= 16'heae5;
assign i[651]= 16'he84c;
assign i[652]= 16'he5b3;
assign i[653]= 16'he329;
assign i[654]= 16'he0b9;
assign i[655]= 16'hde70;
assign i[656]= 16'hdc5b;
assign i[657]= 16'hda83;
assign i[658]= 16'hd8f4;
assign i[659]= 16'hd7b6;
assign i[660]= 16'hd6d2;
assign i[661]= 16'hd64f;
assign i[662]= 16'hd632;
assign i[663]= 16'hd67f;
assign i[664]= 16'hd738;
assign i[665]= 16'hd85d;
assign i[666]= 16'hd9ee;
assign i[667]= 16'hdbe8;
assign i[668]= 16'hde45;
assign i[669]= 16'he0ff;
assign i[670]= 16'he40f;
assign i[671]= 16'he76a;
assign i[672]= 16'heb07;
assign i[673]= 16'heed9;
assign i[674]= 16'hf2d5;
assign i[675]= 16'hf6ed;
assign i[676]= 16'hfb15;
assign i[677]= 16'hff41;
assign i[678]= 16'h363;
assign i[679]= 16'h771;
assign i[680]= 16'hb61;
assign i[681]= 16'hf28;
assign i[682]= 16'h12be;
assign i[683]= 16'h161d;
assign i[684]= 16'h1940;
assign i[685]= 16'h1c23;
assign i[686]= 16'h1ec2;
assign i[687]= 16'h211e;
assign i[688]= 16'h2337;
assign i[689]= 16'h250d;
assign i[690]= 16'h26a4;
assign i[691]= 16'h27ff;
assign i[692]= 16'h2921;
assign i[693]= 16'h2a0f;
assign i[694]= 16'h2acd;
assign i[695]= 16'h2b61;
assign i[696]= 16'h2bcf;
assign i[697]= 16'h2c1c;
assign i[698]= 16'h2c4e;
assign i[699]= 16'h2c69;
assign i[700]= 16'h2c71;
assign i[701]= 16'h2c6c;
assign i[702]= 16'h2c5e;
assign i[703]= 16'h2c4b;
assign i[704]= 16'h2c37;
assign i[705]= 16'h2c25;
assign i[706]= 16'h2c1a;
assign i[707]= 16'h2c19;
assign i[708]= 16'h2c24;
assign i[709]= 16'h2c3e;
assign i[710]= 16'h2c68;
assign i[711]= 16'h2ca4;
assign i[712]= 16'h2cf2;
assign i[713]= 16'h2d51;
assign i[714]= 16'h2dbe;
assign i[715]= 16'h2e38;
assign i[716]= 16'h2eba;
assign i[717]= 16'h2f3f;
assign i[718]= 16'h2fc0;
assign i[719]= 16'h3037;
assign i[720]= 16'h309c;
assign i[721]= 16'h30e6;
assign i[722]= 16'h310c;
assign i[723]= 16'h3108;
assign i[724]= 16'h30d1;
assign i[725]= 16'h305f;
assign i[726]= 16'h2faf;
assign i[727]= 16'h2ebb;
assign i[728]= 16'h2d83;
assign i[729]= 16'h2c07;
assign i[730]= 16'h2a49;
assign i[731]= 16'h2850;
assign i[732]= 16'h2623;
assign i[733]= 16'h23cd;
assign i[734]= 16'h2159;
assign i[735]= 16'h1ed7;
assign i[736]= 16'h1c56;
assign i[737]= 16'h19e6;
assign i[738]= 16'h1796;
assign i[739]= 16'h1577;
assign i[740]= 16'h1397;
assign i[741]= 16'h1202;
assign i[742]= 16'h10c2;
assign i[743]= 16'hfdd;
assign i[744]= 16'hf55;
assign i[745]= 16'hf2a;
assign i[746]= 16'hf56;
assign i[747]= 16'hfcf;
assign i[748]= 16'h1089;
assign i[749]= 16'h1171;
assign i[750]= 16'h1274;
assign i[751]= 16'h137b;
assign i[752]= 16'h146d;
assign i[753]= 16'h1533;
assign i[754]= 16'h15b4;
assign i[755]= 16'h15d9;
assign i[756]= 16'h158d;
assign i[757]= 16'h14bf;
assign i[758]= 16'h1364;
assign i[759]= 16'h1172;
assign i[760]= 16'hee9;
assign i[761]= 16'hbcc;
assign i[762]= 16'h824;
assign i[763]= 16'h403;
assign i[764]= 16'hff7e;
assign i[765]= 16'hfaae;
assign i[766]= 16'hf5b3;
assign i[767]= 16'hf0af;
assign i[768]= 16'hebc7;
assign i[769]= 16'he720;
assign i[770]= 16'he2df;
assign i[771]= 16'hdf27;
assign i[772]= 16'hdc17;
assign i[773]= 16'hd9cd;
assign i[774]= 16'hd85f;
assign i[775]= 16'hd7de;
assign i[776]= 16'hd853;
assign i[777]= 16'hd9c2;
assign i[778]= 16'hdc26;
assign i[779]= 16'hdf73;
assign i[780]= 16'he397;
assign i[781]= 16'he877;
assign i[782]= 16'hedf7;
assign i[783]= 16'hf3f2;
assign i[784]= 16'hfa43;
assign i[785]= 16'hc0;
assign i[786]= 16'h742;
assign i[787]= 16'hda1;
assign i[788]= 16'h13b5;
assign i[789]= 16'h195c;
assign i[790]= 16'h1e75;
assign i[791]= 16'h22e8;
assign i[792]= 16'h26a0;
assign i[793]= 16'h298f;
assign i[794]= 16'h2bac;
assign i[795]= 16'h2cf8;
assign i[796]= 16'h2d76;
assign i[797]= 16'h2d32;
assign i[798]= 16'h2c3b;
assign i[799]= 16'h2aa6;
assign i[800]= 16'h288a;
assign i[801]= 16'h2602;
assign i[802]= 16'h232a;
assign i[803]= 16'h201d;
assign i[804]= 16'h1cf7;
assign i[805]= 16'h19d3;
assign i[806]= 16'h16c9;
assign i[807]= 16'h13ed;
assign i[808]= 16'h1152;
assign i[809]= 16'hf07;
assign i[810]= 16'hd14;
assign i[811]= 16'hb80;
assign i[812]= 16'ha4d;
assign i[813]= 16'h97a;
assign i[814]= 16'h902;
assign i[815]= 16'h8dc;
assign i[816]= 16'h900;
assign i[817]= 16'h95f;
assign i[818]= 16'h9ed;
assign i[819]= 16'ha9c;
assign i[820]= 16'hb5c;
assign i[821]= 16'hc1e;
assign i[822]= 16'hcd5;
assign i[823]= 16'hd73;
assign i[824]= 16'hdec;
assign i[825]= 16'he35;
assign i[826]= 16'he45;
assign i[827]= 16'he15;
assign i[828]= 16'hd9e;
assign i[829]= 16'hcdb;
assign i[830]= 16'hbcb;
assign i[831]= 16'ha6c;
assign i[832]= 16'h8be;
assign i[833]= 16'h6c3;
assign i[834]= 16'h47d;
assign i[835]= 16'h1f2;
assign i[836]= 16'hff27;
assign i[837]= 16'hfc22;
assign i[838]= 16'hf8ec;
assign i[839]= 16'hf58e;
assign i[840]= 16'hf214;
assign i[841]= 16'hee88;
assign i[842]= 16'heaf8;
assign i[843]= 16'he772;
assign i[844]= 16'he404;
assign i[845]= 16'he0bf;
assign i[846]= 16'hddb2;
assign i[847]= 16'hdaed;
assign i[848]= 16'hd881;
assign i[849]= 16'hd67d;
assign i[850]= 16'hd4ef;
assign i[851]= 16'hd3e5;
assign i[852]= 16'hd36a;
assign i[853]= 16'hd388;
assign i[854]= 16'hd446;
assign i[855]= 16'hd5a7;
assign i[856]= 16'hd7ae;
assign i[857]= 16'hda56;
assign i[858]= 16'hdd9c;
assign i[859]= 16'he175;
assign i[860]= 16'he5d6;
assign i[861]= 16'heaaf;
assign i[862]= 16'hefee;
assign i[863]= 16'hf57e;
assign i[864]= 16'hfb49;
assign i[865]= 16'h136;
assign i[866]= 16'h72e;
assign i[867]= 16'hd18;
assign i[868]= 16'h12dc;
assign i[869]= 16'h1862;
assign i[870]= 16'h1d96;
assign i[871]= 16'h2264;
assign i[872]= 16'h26bd;
assign i[873]= 16'h2a94;
assign i[874]= 16'h2de0;
assign i[875]= 16'h309b;
assign i[876]= 16'h32c3;
assign i[877]= 16'h345b;
assign i[878]= 16'h3568;
assign i[879]= 16'h35f3;
assign i[880]= 16'h3607;
assign i[881]= 16'h35b3;
assign i[882]= 16'h3507;
assign i[883]= 16'h3414;
assign i[884]= 16'h32ed;
assign i[885]= 16'h31a3;
assign i[886]= 16'h3048;
assign i[887]= 16'h2eee;
assign i[888]= 16'h2da3;
assign i[889]= 16'h2c74;
assign i[890]= 16'h2b6d;
assign i[891]= 16'h2a96;
assign i[892]= 16'h29f4;
assign i[893]= 16'h2989;
assign i[894]= 16'h2957;
assign i[895]= 16'h2959;
assign i[896]= 16'h298b;
assign i[897]= 16'h29e4;
assign i[898]= 16'h2a5d;
assign i[899]= 16'h2ae9;
assign i[900]= 16'h2b7d;
assign i[901]= 16'h2c0c;
assign i[902]= 16'h2c8a;
assign i[903]= 16'h2ceb;
assign i[904]= 16'h2d23;
assign i[905]= 16'h2d28;
assign i[906]= 16'h2cf1;
assign i[907]= 16'h2c76;
assign i[908]= 16'h2bb1;
assign i[909]= 16'h2aa0;
assign i[910]= 16'h293f;
assign i[911]= 16'h2790;
assign i[912]= 16'h2595;
assign i[913]= 16'h2350;
assign i[914]= 16'h20c7;
assign i[915]= 16'h1e00;
assign i[916]= 16'h1b03;
assign i[917]= 16'h17d6;
assign i[918]= 16'h1483;
assign i[919]= 16'h1110;
assign i[920]= 16'hd86;
assign i[921]= 16'h9ed;
assign i[922]= 16'h64c;
assign i[923]= 16'h2a7;
assign i[924]= 16'hff08;
assign i[925]= 16'hfb6f;
assign i[926]= 16'hf7e3;
assign i[927]= 16'hf466;
assign i[928]= 16'hf0fd;
assign i[929]= 16'heda9;
assign i[930]= 16'hea6e;
assign i[931]= 16'he750;
assign i[932]= 16'he452;
assign i[933]= 16'he177;
assign i[934]= 16'hdec6;
assign i[935]= 16'hdc45;
assign i[936]= 16'hd9fa;
assign i[937]= 16'hd7ee;
assign i[938]= 16'hd62b;
assign i[939]= 16'hd4b9;
assign i[940]= 16'hd3a4;
assign i[941]= 16'hd2f7;
assign i[942]= 16'hd2bd;
assign i[943]= 16'hd2ff;
assign i[944]= 16'hd3c7;
assign i[945]= 16'hd51d;
assign i[946]= 16'hd706;
assign i[947]= 16'hd985;
assign i[948]= 16'hdc9b;
assign i[949]= 16'he043;
assign i[950]= 16'he478;
assign i[951]= 16'he92d;
assign i[952]= 16'hee53;
assign i[953]= 16'hf3d8;
assign i[954]= 16'hf9a4;
assign i[955]= 16'hff9d;
assign i[956]= 16'h5a5;
assign i[957]= 16'hb9e;
assign i[958]= 16'h1167;
assign i[959]= 16'h16dd;
assign i[960]= 16'h1be0;
assign i[961]= 16'h204f;
assign i[962]= 16'h240d;
assign i[963]= 16'h2700;
assign i[964]= 16'h2911;
assign i[965]= 16'h2a31;
assign i[966]= 16'h2a53;
assign i[967]= 16'h2974;
assign i[968]= 16'h2796;
assign i[969]= 16'h24c2;
assign i[970]= 16'h2109;
assign i[971]= 16'h1c81;
assign i[972]= 16'h1748;
assign i[973]= 16'h117f;
assign i[974]= 16'hb4f;
assign i[975]= 16'h4e1;
assign i[976]= 16'hfe63;
assign i[977]= 16'hf801;
assign i[978]= 16'hf1e9;
assign i[979]= 16'hec47;
assign i[980]= 16'he743;
assign i[981]= 16'he301;
assign i[982]= 16'hdfa2;
assign i[983]= 16'hdd3c;
assign i[984]= 16'hdbe1;
assign i[985]= 16'hdb9c;
assign i[986]= 16'hdc6e;
assign i[987]= 16'hde53;
assign i[988]= 16'he13b;
assign i[989]= 16'he514;
assign i[990]= 16'he9c2;
assign i[991]= 16'hef25;
assign i[992]= 16'hf518;
assign i[993]= 16'hfb72;
assign i[994]= 16'h20a;
assign i[995]= 16'h8b5;
assign i[996]= 16'hf48;
assign i[997]= 16'h159c;
assign i[998]= 16'h1b89;
assign i[999]= 16'h20ef;
assign i[1000]= 16'h25b0;
assign i[1001]= 16'h29b4;
assign i[1002]= 16'h2ceb;
assign i[1003]= 16'h2f47;
assign i[1004]= 16'h30c4;
assign i[1005]= 16'h3163;
assign i[1006]= 16'h3128;
assign i[1007]= 16'h3020;
assign i[1008]= 16'h2e5a;
assign i[1009]= 16'h2bea;
assign i[1010]= 16'h28e7;
assign i[1011]= 16'h2568;
assign i[1012]= 16'h2189;
assign i[1013]= 16'h1d64;
assign i[1014]= 16'h1912;
assign i[1015]= 16'h14ad;
assign i[1016]= 16'h104e;
assign i[1017]= 16'hc09;
assign i[1018]= 16'h7f3;
assign i[1019]= 16'h41b;
assign i[1020]= 16'h90;
assign i[1021]= 16'hfd5e;
assign i[1022]= 16'hfa8c;
assign i[1023]= 16'hf821;
assign i[1024]= 16'hf620;
assign i[1025]= 16'hf48b;
assign i[1026]= 16'hf361;
assign i[1027]= 16'hf2a0;
assign i[1028]= 16'hf245;
assign i[1029]= 16'hf24a;
assign i[1030]= 16'hf2aa;
assign i[1031]= 16'hf35e;
assign i[1032]= 16'hf45d;
assign i[1033]= 16'hf5a1;
assign i[1034]= 16'hf71e;
assign i[1035]= 16'hf8cd;
assign i[1036]= 16'hfaa1;
assign i[1037]= 16'hfc90;
assign i[1038]= 16'hfe8f;
assign i[1039]= 16'h91;
assign i[1040]= 16'h28b;
assign i[1041]= 16'h46f;
assign i[1042]= 16'h632;
assign i[1043]= 16'h7c8;
assign i[1044]= 16'h924;
assign i[1045]= 16'ha3d;
assign i[1046]= 16'hb0a;
assign i[1047]= 16'hb84;
assign i[1048]= 16'hba4;
assign i[1049]= 16'hb6a;
assign i[1050]= 16'had3;
assign i[1051]= 16'h9e3;
assign i[1052]= 16'h89f;
assign i[1053]= 16'h710;
assign i[1054]= 16'h540;
assign i[1055]= 16'h33e;
assign i[1056]= 16'h118;
assign i[1057]= 16'hfee2;
assign i[1058]= 16'hfcad;
assign i[1059]= 16'hfa8c;
assign i[1060]= 16'hf892;
assign i[1061]= 16'hf6d4;
assign i[1062]= 16'hf560;
assign i[1063]= 16'hf446;
assign i[1064]= 16'hf392;
assign i[1065]= 16'hf34d;
assign i[1066]= 16'hf37a;
assign i[1067]= 16'hf41a;
assign i[1068]= 16'hf52b;
assign i[1069]= 16'hf6a3;
assign i[1070]= 16'hf877;
assign i[1071]= 16'hfa97;
assign i[1072]= 16'hfcf2;
assign i[1073]= 16'hff71;
assign i[1074]= 16'h1fd;
assign i[1075]= 16'h47f;
assign i[1076]= 16'h6e0;
assign i[1077]= 16'h907;
assign i[1078]= 16'hae1;
assign i[1079]= 16'hc5b;
assign i[1080]= 16'hd66;
assign i[1081]= 16'hdf6;
assign i[1082]= 16'he05;
assign i[1083]= 16'hd92;
assign i[1084]= 16'hc9f;
assign i[1085]= 16'hb33;
assign i[1086]= 16'h95b;
assign i[1087]= 16'h726;
assign i[1088]= 16'h4a8;
assign i[1089]= 16'h1f6;
assign i[1090]= 16'hff27;
assign i[1091]= 16'hfc52;
assign i[1092]= 16'hf98e;
assign i[1093]= 16'hf6f2;
assign i[1094]= 16'hf492;
assign i[1095]= 16'hf27d;
assign i[1096]= 16'hf0c0;
assign i[1097]= 16'hef65;
assign i[1098]= 16'hee70;
assign i[1099]= 16'hede0;
assign i[1100]= 16'hedb1;
assign i[1101]= 16'hedd8;
assign i[1102]= 16'hee4a;
assign i[1103]= 16'heef7;
assign i[1104]= 16'hefcb;
assign i[1105]= 16'hf0b3;
assign i[1106]= 16'hf19c;
assign i[1107]= 16'hf272;
assign i[1108]= 16'hf323;
assign i[1109]= 16'hf3a0;
assign i[1110]= 16'hf3dc;
assign i[1111]= 16'hf3cf;
assign i[1112]= 16'hf377;
assign i[1113]= 16'hf2d3;
assign i[1114]= 16'hf1ea;
assign i[1115]= 16'hf0c6;
assign i[1116]= 16'hef75;
assign i[1117]= 16'hee0c;
assign i[1118]= 16'hec9f;
assign i[1119]= 16'heb46;
assign i[1120]= 16'hea19;
assign i[1121]= 16'he933;
assign i[1122]= 16'he8a9;
assign i[1123]= 16'he892;
assign i[1124]= 16'he901;
assign i[1125]= 16'hea02;
assign i[1126]= 16'heba0;
assign i[1127]= 16'heddd;
assign i[1128]= 16'hf0b8;
assign i[1129]= 16'hf428;
assign i[1130]= 16'hf81f;
assign i[1131]= 16'hfc89;
assign i[1132]= 16'h14b;
assign i[1133]= 16'h64a;
assign i[1134]= 16'hb64;
assign i[1135]= 16'h1075;
assign i[1136]= 16'h1559;
assign i[1137]= 16'h19eb;
assign i[1138]= 16'h1e08;
assign i[1139]= 16'h218e;
assign i[1140]= 16'h2461;
assign i[1141]= 16'h2667;
assign i[1142]= 16'h278f;
assign i[1143]= 16'h27cb;
assign i[1144]= 16'h2714;
assign i[1145]= 16'h256c;
assign i[1146]= 16'h22da;
assign i[1147]= 16'h1f6d;
assign i[1148]= 16'h1b38;
assign i[1149]= 16'h1655;
assign i[1150]= 16'h10e4;
assign i[1151]= 16'hb08;
assign i[1152]= 16'h4e4;
assign i[1153]= 16'hfea2;
assign i[1154]= 16'hf866;
assign i[1155]= 16'hf258;
assign i[1156]= 16'hec9e;
assign i[1157]= 16'he759;
assign i[1158]= 16'he2a9;
assign i[1159]= 16'hdea8;
assign i[1160]= 16'hdb6b;
assign i[1161]= 16'hd903;
assign i[1162]= 16'hd77b;
assign i[1163]= 16'hd6d8;
assign i[1164]= 16'hd71b;
assign i[1165]= 16'hd83e;
assign i[1166]= 16'hda38;
assign i[1167]= 16'hdcfb;
assign i[1168]= 16'he076;
assign i[1169]= 16'he493;
assign i[1170]= 16'he93c;
assign i[1171]= 16'hee57;
assign i[1172]= 16'hf3cc;
assign i[1173]= 16'hf97f;
assign i[1174]= 16'hff56;
assign i[1175]= 16'h536;
assign i[1176]= 16'hb08;
assign i[1177]= 16'h10b2;
assign i[1178]= 16'h161f;
assign i[1179]= 16'h1b39;
assign i[1180]= 16'h1fed;
assign i[1181]= 16'h2429;
assign i[1182]= 16'h27df;
assign i[1183]= 16'h2b01;
assign i[1184]= 16'h2d84;
assign i[1185]= 16'h2f5e;
assign i[1186]= 16'h3089;
assign i[1187]= 16'h3100;
assign i[1188]= 16'h30c0;
assign i[1189]= 16'h2fca;
assign i[1190]= 16'h2e1f;
assign i[1191]= 16'h2bc5;
assign i[1192]= 16'h28c4;
assign i[1193]= 16'h2525;
assign i[1194]= 16'h20f6;
assign i[1195]= 16'h1c46;
assign i[1196]= 16'h1728;
assign i[1197]= 16'h11af;
assign i[1198]= 16'hbf4;
assign i[1199]= 16'h60d;
assign i[1200]= 16'h14;
assign i[1201]= 16'hfa24;
assign i[1202]= 16'hf457;
assign i[1203]= 16'heec6;
assign i[1204]= 16'he98c;
assign i[1205]= 16'he4be;
assign i[1206]= 16'he073;
assign i[1207]= 16'hdcbb;
assign i[1208]= 16'hd9a5;
assign i[1209]= 16'hd73c;
assign i[1210]= 16'hd586;
assign i[1211]= 16'hd485;
assign i[1212]= 16'hd435;
assign i[1213]= 16'hd48f;
assign i[1214]= 16'hd589;
assign i[1215]= 16'hd713;
assign i[1216]= 16'hd91a;
assign i[1217]= 16'hdb8b;
assign i[1218]= 16'hde4d;
assign i[1219]= 16'he14b;
assign i[1220]= 16'he46c;
assign i[1221]= 16'he79a;
assign i[1222]= 16'heabf;
assign i[1223]= 16'hedc9;
assign i[1224]= 16'hf0a8;
assign i[1225]= 16'hf350;
assign i[1226]= 16'hf5ba;
assign i[1227]= 16'hf7e2;
assign i[1228]= 16'hf9c8;
assign i[1229]= 16'hfb71;
assign i[1230]= 16'hfce4;
assign i[1231]= 16'hfe2f;
assign i[1232]= 16'hff5e;
assign i[1233]= 16'h81;
assign i[1234]= 16'h1aa;
assign i[1235]= 16'h2e9;
assign i[1236]= 16'h44d;
assign i[1237]= 16'h5e3;
assign i[1238]= 16'h7b8;
assign i[1239]= 16'h9d1;
assign i[1240]= 16'hc33;
assign i[1241]= 16'hedc;
assign i[1242]= 16'h11c6;
assign i[1243]= 16'h14e6;
assign i[1244]= 16'h182f;
assign i[1245]= 16'h1b8c;
assign i[1246]= 16'h1ee7;
assign i[1247]= 16'h2227;
assign i[1248]= 16'h2530;
assign i[1249]= 16'h27e8;
assign i[1250]= 16'h2a33;
assign i[1251]= 16'h2bf7;
assign i[1252]= 16'h2d1c;
assign i[1253]= 16'h2d8e;
assign i[1254]= 16'h2d3f;
assign i[1255]= 16'h2c23;
assign i[1256]= 16'h2a36;
assign i[1257]= 16'h277a;
assign i[1258]= 16'h23f5;
assign i[1259]= 16'h1fb6;
assign i[1260]= 16'h1acf;
assign i[1261]= 16'h1559;
assign i[1262]= 16'hf71;
assign i[1263]= 16'h937;
assign i[1264]= 16'h2ce;
assign i[1265]= 16'hfc5a;
assign i[1266]= 16'hf600;
assign i[1267]= 16'hefe2;
assign i[1268]= 16'hea22;
assign i[1269]= 16'he4de;
assign i[1270]= 16'he031;
assign i[1271]= 16'hdc2f;
assign i[1272]= 16'hd8e9;
assign i[1273]= 16'hd668;
assign i[1274]= 16'hd4b0;
assign i[1275]= 16'hd3c1;
assign i[1276]= 16'hd391;
assign i[1277]= 16'hd416;
assign i[1278]= 16'hd53e;
assign i[1279]= 16'hd6f4;
assign i[1280]= 16'hd91f;
assign i[1281]= 16'hdba7;
assign i[1282]= 16'hde70;
assign i[1283]= 16'he160;
assign i[1284]= 16'he45b;
assign i[1285]= 16'he749;
assign i[1286]= 16'hea15;
assign i[1287]= 16'hecac;
assign i[1288]= 16'heefc;
assign i[1289]= 16'hf0fc;
assign i[1290]= 16'hf2a3;
assign i[1291]= 16'hf3ee;
assign i[1292]= 16'hf4dc;
assign i[1293]= 16'hf572;
assign i[1294]= 16'hf5b6;
assign i[1295]= 16'hf5b3;
assign i[1296]= 16'hf573;
assign i[1297]= 16'hf506;
assign i[1298]= 16'hf479;
assign i[1299]= 16'hf3db;
assign i[1300]= 16'hf33c;
assign i[1301]= 16'hf2a9;
assign i[1302]= 16'hf230;
assign i[1303]= 16'hf1dc;
assign i[1304]= 16'hf1b8;
assign i[1305]= 16'hf1cb;
assign i[1306]= 16'hf21d;
assign i[1307]= 16'hf2b0;
assign i[1308]= 16'hf388;
assign i[1309]= 16'hf4a5;
assign i[1310]= 16'hf605;
assign i[1311]= 16'hf7a6;
assign i[1312]= 16'hf984;
assign i[1313]= 16'hfb99;
assign i[1314]= 16'hfde0;
assign i[1315]= 16'h52;
assign i[1316]= 16'h2ea;
assign i[1317]= 16'h59f;
assign i[1318]= 16'h86a;
assign i[1319]= 16'hb44;
assign i[1320]= 16'he25;
assign i[1321]= 16'h1107;
assign i[1322]= 16'h13e1;
assign i[1323]= 16'h16ad;
assign i[1324]= 16'h1963;
assign i[1325]= 16'h1bfc;
assign i[1326]= 16'h1e72;
assign i[1327]= 16'h20be;
assign i[1328]= 16'h22d9;
assign i[1329]= 16'h24bc;
assign i[1330]= 16'h2663;
assign i[1331]= 16'h27c7;
assign i[1332]= 16'h28e5;
assign i[1333]= 16'h29b8;
assign i[1334]= 16'h2a3d;
assign i[1335]= 16'h2a74;
assign i[1336]= 16'h2a5c;
assign i[1337]= 16'h29f6;
assign i[1338]= 16'h2944;
assign i[1339]= 16'h284b;
assign i[1340]= 16'h2711;
assign i[1341]= 16'h259b;
assign i[1342]= 16'h23f2;
assign i[1343]= 16'h2220;
assign i[1344]= 16'h202f;
assign i[1345]= 16'h1e2a;
assign i[1346]= 16'h1c1b;
assign i[1347]= 16'h1a0f;
assign i[1348]= 16'h1810;
assign i[1349]= 16'h1628;
assign i[1350]= 16'h1460;
assign i[1351]= 16'h12c2;
assign i[1352]= 16'h1152;
assign i[1353]= 16'h1017;
assign i[1354]= 16'hf12;
assign i[1355]= 16'he45;
assign i[1356]= 16'hdb0;
assign i[1357]= 16'hd4f;
assign i[1358]= 16'hd1d;
assign i[1359]= 16'hd14;
assign i[1360]= 16'hd2c;
assign i[1361]= 16'hd5d;
assign i[1362]= 16'hd9d;
assign i[1363]= 16'hde2;
assign i[1364]= 16'he21;
assign i[1365]= 16'he50;
assign i[1366]= 16'he65;
assign i[1367]= 16'he59;
assign i[1368]= 16'he22;
assign i[1369]= 16'hdbc;
assign i[1370]= 16'hd21;
assign i[1371]= 16'hc4d;
assign i[1372]= 16'hb40;
assign i[1373]= 16'h9f8;
assign i[1374]= 16'h878;
assign i[1375]= 16'h6c2;
assign i[1376]= 16'h4db;
assign i[1377]= 16'h2c7;
assign i[1378]= 16'h8e;
assign i[1379]= 16'hfe36;
assign i[1380]= 16'hfbc5;
assign i[1381]= 16'hf943;
assign i[1382]= 16'hf6b7;
assign i[1383]= 16'hf427;
assign i[1384]= 16'hf19c;
assign i[1385]= 16'hef1a;
assign i[1386]= 16'heca6;
assign i[1387]= 16'hea45;
assign i[1388]= 16'he7fa;
assign i[1389]= 16'he5c9;
assign i[1390]= 16'he3b4;
assign i[1391]= 16'he1bb;
assign i[1392]= 16'hdfe0;
assign i[1393]= 16'hde22;
assign i[1394]= 16'hdc83;
assign i[1395]= 16'hdb01;
assign i[1396]= 16'hd99c;
assign i[1397]= 16'hd854;
assign i[1398]= 16'hd727;
assign i[1399]= 16'hd615;
assign i[1400]= 16'hd51d;
assign i[1401]= 16'hd440;
assign i[1402]= 16'hd37c;
assign i[1403]= 16'hd2d2;
assign i[1404]= 16'hd241;
assign i[1405]= 16'hd1c9;
assign i[1406]= 16'hd169;
assign i[1407]= 16'hd122;
assign i[1408]= 16'hd0f3;
assign i[1409]= 16'hd0da;
assign i[1410]= 16'hd0d8;
assign i[1411]= 16'hd0e9;
assign i[1412]= 16'hd10d;
assign i[1413]= 16'hd141;
assign i[1414]= 16'hd183;
assign i[1415]= 16'hd1cf;
assign i[1416]= 16'hd224;
assign i[1417]= 16'hd27c;
assign i[1418]= 16'hd2d5;
assign i[1419]= 16'hd32c;
assign i[1420]= 16'hd37d;
assign i[1421]= 16'hd3c5;
assign i[1422]= 16'hd401;
assign i[1423]= 16'hd42f;
assign i[1424]= 16'hd44c;
assign i[1425]= 16'hd458;
assign i[1426]= 16'hd451;
assign i[1427]= 16'hd438;
assign i[1428]= 16'hd40c;
assign i[1429]= 16'hd3d0;
assign i[1430]= 16'hd384;
assign i[1431]= 16'hd32c;
assign i[1432]= 16'hd2ca;
assign i[1433]= 16'hd262;
assign i[1434]= 16'hd1f8;
assign i[1435]= 16'hd190;
assign i[1436]= 16'hd12e;
assign i[1437]= 16'hd0d7;
assign i[1438]= 16'hd090;
assign i[1439]= 16'hd05b;
assign i[1440]= 16'hd03f;
assign i[1441]= 16'hd03d;
assign i[1442]= 16'hd059;
assign i[1443]= 16'hd097;
assign i[1444]= 16'hd0f8;
assign i[1445]= 16'hd17d;
assign i[1446]= 16'hd229;
assign i[1447]= 16'hd2fa;
assign i[1448]= 16'hd3f1;
assign i[1449]= 16'hd50c;
assign i[1450]= 16'hd64b;
assign i[1451]= 16'hd7ab;
assign i[1452]= 16'hd928;
assign i[1453]= 16'hdac2;
assign i[1454]= 16'hdc72;
assign i[1455]= 16'hde37;
assign i[1456]= 16'he00a;
assign i[1457]= 16'he1e8;
assign i[1458]= 16'he3cc;
assign i[1459]= 16'he5b0;
assign i[1460]= 16'he791;
assign i[1461]= 16'he967;
assign i[1462]= 16'heb2f;
assign i[1463]= 16'hece2;
assign i[1464]= 16'hee7d;
assign i[1465]= 16'heffa;
assign i[1466]= 16'hf154;
assign i[1467]= 16'hf287;
assign i[1468]= 16'hf38f;
assign i[1469]= 16'hf469;
assign i[1470]= 16'hf511;
assign i[1471]= 16'hf585;
assign i[1472]= 16'hf5c3;
assign i[1473]= 16'hf5cb;
assign i[1474]= 16'hf59b;
assign i[1475]= 16'hf534;
assign i[1476]= 16'hf496;
assign i[1477]= 16'hf3c4;
assign i[1478]= 16'hf2c1;
assign i[1479]= 16'hf18f;
assign i[1480]= 16'hf032;
assign i[1481]= 16'heeaf;
assign i[1482]= 16'hed0c;
assign i[1483]= 16'heb4d;
assign i[1484]= 16'he978;
assign i[1485]= 16'he794;
assign i[1486]= 16'he5a6;
assign i[1487]= 16'he3b6;
assign i[1488]= 16'he1c8;
assign i[1489]= 16'hdfe2;
assign i[1490]= 16'hde0a;
assign i[1491]= 16'hdc45;
assign i[1492]= 16'hda97;
assign i[1493]= 16'hd903;
assign i[1494]= 16'hd78e;
assign i[1495]= 16'hd638;
assign i[1496]= 16'hd504;
assign i[1497]= 16'hd3f3;
assign i[1498]= 16'hd306;
assign i[1499]= 16'hd23c;
assign i[1500]= 16'hd195;
assign i[1501]= 16'hd110;
assign i[1502]= 16'hd0ab;
assign i[1503]= 16'hd066;
assign i[1504]= 16'hd03d;
assign i[1505]= 16'hd02f;
assign i[1506]= 16'hd03a;
assign i[1507]= 16'hd05c;
assign i[1508]= 16'hd092;
assign i[1509]= 16'hd0d9;
assign i[1510]= 16'hd12f;
assign i[1511]= 16'hd192;
assign i[1512]= 16'hd1fe;
assign i[1513]= 16'hd271;
assign i[1514]= 16'hd2e7;
assign i[1515]= 16'hd35d;
assign i[1516]= 16'hd3d0;
assign i[1517]= 16'hd43d;
assign i[1518]= 16'hd49e;
assign i[1519]= 16'hd4f1;
assign i[1520]= 16'hd532;
assign i[1521]= 16'hd55d;
assign i[1522]= 16'hd56f;
assign i[1523]= 16'hd566;
assign i[1524]= 16'hd53f;
assign i[1525]= 16'hd4f9;
assign i[1526]= 16'hd494;
assign i[1527]= 16'hd412;
assign i[1528]= 16'hd373;
assign i[1529]= 16'hd2bc;
assign i[1530]= 16'hd1f2;
assign i[1531]= 16'hd11b;
assign i[1532]= 16'hd040;
assign i[1533]= 16'hcf69;
assign i[1534]= 16'hcea2;
assign i[1535]= 16'hcdf5;
assign i[1536]= 16'hcd6e;
assign i[1537]= 16'hcd1a;
assign i[1538]= 16'hcd03;
assign i[1539]= 16'hcd36;
assign i[1540]= 16'hcdbd;
assign i[1541]= 16'hcea0;
assign i[1542]= 16'hcfe6;
assign i[1543]= 16'hd193;
assign i[1544]= 16'hd3aa;
assign i[1545]= 16'hd629;
assign i[1546]= 16'hd90c;
assign i[1547]= 16'hdc4c;
assign i[1548]= 16'hdfe0;
assign i[1549]= 16'he3bb;
assign i[1550]= 16'he7cc;
assign i[1551]= 16'hec04;
assign i[1552]= 16'hf04e;
assign i[1553]= 16'hf497;
assign i[1554]= 16'hf8cb;
assign i[1555]= 16'hfcd6;
assign i[1556]= 16'ha3;
assign i[1557]= 16'h424;
assign i[1558]= 16'h749;
assign i[1559]= 16'ha06;
assign i[1560]= 16'hc53;
assign i[1561]= 16'he2b;
assign i[1562]= 16'hf8d;
assign i[1563]= 16'h107e;
assign i[1564]= 16'h1104;
assign i[1565]= 16'h112b;
assign i[1566]= 16'h1102;
assign i[1567]= 16'h1099;
assign i[1568]= 16'h1005;
assign i[1569]= 16'hf5a;
assign i[1570]= 16'heae;
assign i[1571]= 16'he15;
assign i[1572]= 16'hda4;
assign i[1573]= 16'hd6e;
assign i[1574]= 16'hd7f;
assign i[1575]= 16'hde6;
assign i[1576]= 16'hea8;
assign i[1577]= 16'hfca;
assign i[1578]= 16'h114a;
assign i[1579]= 16'h1323;
assign i[1580]= 16'h154a;
assign i[1581]= 16'h17b2;
assign i[1582]= 16'h1a49;
assign i[1583]= 16'h1cfa;
assign i[1584]= 16'h1fb0;
assign i[1585]= 16'h2254;
assign i[1586]= 16'h24ce;
assign i[1587]= 16'h2707;
assign i[1588]= 16'h28ec;
assign i[1589]= 16'h2a6a;
assign i[1590]= 16'h2b74;
assign i[1591]= 16'h2bff;
assign i[1592]= 16'h2c06;
assign i[1593]= 16'h2b89;
assign i[1594]= 16'h2a8b;
assign i[1595]= 16'h2917;
assign i[1596]= 16'h273b;
assign i[1597]= 16'h2509;
assign i[1598]= 16'h2297;
assign i[1599]= 16'h1ffc;
assign i[1600]= 16'h1d53;
assign i[1601]= 16'h1ab6;
assign i[1602]= 16'h183f;
assign i[1603]= 16'h1608;
assign i[1604]= 16'h1425;
assign i[1605]= 16'h12aa;
assign i[1606]= 16'h11a6;
assign i[1607]= 16'h1124;
assign i[1608]= 16'h1127;
assign i[1609]= 16'h11af;
assign i[1610]= 16'h12b8;
assign i[1611]= 16'h1435;
assign i[1612]= 16'h1618;
assign i[1613]= 16'h184d;
assign i[1614]= 16'h1abb;
assign i[1615]= 16'h1d48;
assign i[1616]= 16'h1fd9;
assign i[1617]= 16'h2251;
assign i[1618]= 16'h2491;
assign i[1619]= 16'h2680;
assign i[1620]= 16'h2803;
assign i[1621]= 16'h2903;
assign i[1622]= 16'h296d;
assign i[1623]= 16'h2933;
assign i[1624]= 16'h2849;
assign i[1625]= 16'h26a9;
assign i[1626]= 16'h2454;
assign i[1627]= 16'h214d;
assign i[1628]= 16'h1d9c;
assign i[1629]= 16'h194f;
assign i[1630]= 16'h1476;
assign i[1631]= 16'hf24;
assign i[1632]= 16'h970;
assign i[1633]= 16'h371;
assign i[1634]= 16'hfd43;
assign i[1635]= 16'hf6fd;
assign i[1636]= 16'hf0b9;
assign i[1637]= 16'hea91;
assign i[1638]= 16'he49c;
assign i[1639]= 16'hdef0;
assign i[1640]= 16'hd9a3;
assign i[1641]= 16'hd4c5;
assign i[1642]= 16'hd067;
assign i[1643]= 16'hcc96;
assign i[1644]= 16'hc95d;
assign i[1645]= 16'hc6c3;
assign i[1646]= 16'hc4ce;
assign i[1647]= 16'hc383;
assign i[1648]= 16'hc2e1;
assign i[1649]= 16'hc2e8;
assign i[1650]= 16'hc395;
assign i[1651]= 16'hc4e2;
assign i[1652]= 16'hc6c8;
assign i[1653]= 16'hc93e;
assign i[1654]= 16'hcc39;
assign i[1655]= 16'hcfac;
assign i[1656]= 16'hd389;
assign i[1657]= 16'hd7bd;
assign i[1658]= 16'hdc39;
assign i[1659]= 16'he0e7;
assign i[1660]= 16'he5b4;
assign i[1661]= 16'hea88;
assign i[1662]= 16'hef4d;
assign i[1663]= 16'hf3ec;
assign i[1664]= 16'hf84e;
assign i[1665]= 16'hfc5c;
assign i[1666]= 16'h0;
assign i[1667]= 16'h326;
assign i[1668]= 16'h5bd;
assign i[1669]= 16'h7b7;
assign i[1670]= 16'h906;
assign i[1671]= 16'h9a4;
assign i[1672]= 16'h98c;
assign i[1673]= 16'h8bf;
assign i[1674]= 16'h742;
assign i[1675]= 16'h520;
assign i[1676]= 16'h267;
assign i[1677]= 16'hff2a;
assign i[1678]= 16'hfb7e;
assign i[1679]= 16'hf77e;
assign i[1680]= 16'hf346;
assign i[1681]= 16'heef3;
assign i[1682]= 16'heaa5;
assign i[1683]= 16'he67a;
assign i[1684]= 16'he28f;
assign i[1685]= 16'hdeff;
assign i[1686]= 16'hdbe3;
assign i[1687]= 16'hd94f;
assign i[1688]= 16'hd753;
assign i[1689]= 16'hd5f9;
assign i[1690]= 16'hd547;
assign i[1691]= 16'hd53a;
assign i[1692]= 16'hd5ce;
assign i[1693]= 16'hd6f6;
assign i[1694]= 16'hd8a1;
assign i[1695]= 16'hdab9;
assign i[1696]= 16'hdd26;
assign i[1697]= 16'hdfcc;
assign i[1698]= 16'he28c;
assign i[1699]= 16'he548;
assign i[1700]= 16'he7e4;
assign i[1701]= 16'hea42;
assign i[1702]= 16'hec49;
assign i[1703]= 16'hede5;
assign i[1704]= 16'hef03;
assign i[1705]= 16'hef98;
assign i[1706]= 16'hef9d;
assign i[1707]= 16'hef12;
assign i[1708]= 16'hedfc;
assign i[1709]= 16'hec65;
assign i[1710]= 16'hea5f;
assign i[1711]= 16'he7fe;
assign i[1712]= 16'he55a;
assign i[1713]= 16'he28d;
assign i[1714]= 16'hdfb6;
assign i[1715]= 16'hdcf0;
assign i[1716]= 16'hda58;
assign i[1717]= 16'hd80a;
assign i[1718]= 16'hd61c;
assign i[1719]= 16'hd4a2;
assign i[1720]= 16'hd3ad;
assign i[1721]= 16'hd345;
assign i[1722]= 16'hd370;
assign i[1723]= 16'hd42b;
assign i[1724]= 16'hd571;
assign i[1725]= 16'hd733;
assign i[1726]= 16'hd962;
assign i[1727]= 16'hdbe8;
assign i[1728]= 16'hdeac;
assign i[1729]= 16'he194;
assign i[1730]= 16'he483;
assign i[1731]= 16'he760;
assign i[1732]= 16'hea0e;
assign i[1733]= 16'hec78;
assign i[1734]= 16'hee89;
assign i[1735]= 16'hf032;
assign i[1736]= 16'hf169;
assign i[1737]= 16'hf228;
assign i[1738]= 16'hf271;
assign i[1739]= 16'hf24c;
assign i[1740]= 16'hf1c5;
assign i[1741]= 16'hf0ee;
assign i[1742]= 16'hefde;
assign i[1743]= 16'heeb0;
assign i[1744]= 16'hed7e;
assign i[1745]= 16'hec69;
assign i[1746]= 16'heb8c;
assign i[1747]= 16'heb05;
assign i[1748]= 16'heaed;
assign i[1749]= 16'heb5b;
assign i[1750]= 16'hec5f;
assign i[1751]= 16'hee05;
assign i[1752]= 16'hf051;
assign i[1753]= 16'hf343;
assign i[1754]= 16'hf6cf;
assign i[1755]= 16'hfae8;
assign i[1756]= 16'hff76;
assign i[1757]= 16'h45d;
assign i[1758]= 16'h97c;
assign i[1759]= 16'heaf;
assign i[1760]= 16'h13cd;
assign i[1761]= 16'h18ae;
assign i[1762]= 16'h1d29;
assign i[1763]= 16'h2119;
assign i[1764]= 16'h245a;
assign i[1765]= 16'h26cc;
assign i[1766]= 16'h2857;
assign i[1767]= 16'h28e9;
assign i[1768]= 16'h2877;
assign i[1769]= 16'h26fd;
assign i[1770]= 16'h2481;
assign i[1771]= 16'h210f;
assign i[1772]= 16'h1cbd;
assign i[1773]= 16'h17a5;
assign i[1774]= 16'h11e9;
assign i[1775]= 16'hbaf;
assign i[1776]= 16'h521;
assign i[1777]= 16'hfe6b;
assign i[1778]= 16'hf7b8;
assign i[1779]= 16'hf135;
assign i[1780]= 16'heb0a;
assign i[1781]= 16'he55c;
assign i[1782]= 16'he04d;
assign i[1783]= 16'hdbf6;
assign i[1784]= 16'hd86c;
assign i[1785]= 16'hd5bc;
assign i[1786]= 16'hd3eb;
assign i[1787]= 16'hd2f8;
assign i[1788]= 16'hd2da;
assign i[1789]= 16'hd381;
assign i[1790]= 16'hd4da;
assign i[1791]= 16'hd6cb;
assign i[1792]= 16'hd938;
assign i[1793]= 16'hdc01;
assign i[1794]= 16'hdf06;
assign i[1795]= 16'he228;
assign i[1796]= 16'he548;
assign i[1797]= 16'he84a;
assign i[1798]= 16'heb15;
assign i[1799]= 16'hed97;
assign i[1800]= 16'hefbe;
assign i[1801]= 16'hf180;
assign i[1802]= 16'hf2da;
assign i[1803]= 16'hf3ca;
assign i[1804]= 16'hf455;
assign i[1805]= 16'hf485;
assign i[1806]= 16'hf467;
assign i[1807]= 16'hf40a;
assign i[1808]= 16'hf381;
assign i[1809]= 16'hf2de;
assign i[1810]= 16'hf236;
assign i[1811]= 16'hf19b;
assign i[1812]= 16'hf11f;
assign i[1813]= 16'hf0d0;
assign i[1814]= 16'hf0bc;
assign i[1815]= 16'hf0eb;
assign i[1816]= 16'hf165;
assign i[1817]= 16'hf22c;
assign i[1818]= 16'hf33f;
assign i[1819]= 16'hf499;
assign i[1820]= 16'hf634;
assign i[1821]= 16'hf806;
assign i[1822]= 16'hfa04;
assign i[1823]= 16'hfc1f;
assign i[1824]= 16'hfe4a;
assign i[1825]= 16'h76;
assign i[1826]= 16'h295;
assign i[1827]= 16'h499;
assign i[1828]= 16'h675;
assign i[1829]= 16'h81e;
assign i[1830]= 16'h989;
assign i[1831]= 16'hab0;
assign i[1832]= 16'hb8c;
assign i[1833]= 16'hc18;
assign i[1834]= 16'hc53;
assign i[1835]= 16'hc3c;
assign i[1836]= 16'hbd3;
assign i[1837]= 16'hb1b;
assign i[1838]= 16'ha16;
assign i[1839]= 16'h8c9;
assign i[1840]= 16'h739;
assign i[1841]= 16'h56c;
assign i[1842]= 16'h368;
assign i[1843]= 16'h134;
assign i[1844]= 16'hfed8;
assign i[1845]= 16'hfc5c;
assign i[1846]= 16'hf9c9;
assign i[1847]= 16'hf729;
assign i[1848]= 16'hf487;
assign i[1849]= 16'hf1ee;
assign i[1850]= 16'hef6b;
assign i[1851]= 16'hed0b;
assign i[1852]= 16'headc;
assign i[1853]= 16'he8ec;
assign i[1854]= 16'he74a;
assign i[1855]= 16'he605;
assign i[1856]= 16'he529;
assign i[1857]= 16'he4c4;
assign i[1858]= 16'he4e1;
assign i[1859]= 16'he588;
assign i[1860]= 16'he6c0;
assign i[1861]= 16'he88c;
assign i[1862]= 16'heaeb;
assign i[1863]= 16'hedd9;
assign i[1864]= 16'hf14e;
assign i[1865]= 16'hf53d;
assign i[1866]= 16'hf994;
assign i[1867]= 16'hfe41;
assign i[1868]= 16'h328;
assign i[1869]= 16'h830;
assign i[1870]= 16'hd3b;
assign i[1871]= 16'h122a;
assign i[1872]= 16'h16dc;
assign i[1873]= 16'h1b31;
assign i[1874]= 16'h1f0c;
assign i[1875]= 16'h224e;
assign i[1876]= 16'h24e0;
assign i[1877]= 16'h26ac;
assign i[1878]= 16'h27a1;
assign i[1879]= 16'h27b5;
assign i[1880]= 16'h26e2;
assign i[1881]= 16'h252a;
assign i[1882]= 16'h2294;
assign i[1883]= 16'h1f2c;
assign i[1884]= 16'h1b05;
assign i[1885]= 16'h1638;
assign i[1886]= 16'h10e0;
assign i[1887]= 16'hb1c;
assign i[1888]= 16'h510;
assign i[1889]= 16'hfedf;
assign i[1890]= 16'hf8ab;
assign i[1891]= 16'hf29a;
assign i[1892]= 16'heccb;
assign i[1893]= 16'he75f;
assign i[1894]= 16'he271;
assign i[1895]= 16'hde17;
assign i[1896]= 16'hda64;
assign i[1897]= 16'hd766;
assign i[1898]= 16'hd524;
assign i[1899]= 16'hd3a2;
assign i[1900]= 16'hd2de;
assign i[1901]= 16'hd2cf;
assign i[1902]= 16'hd36c;
assign i[1903]= 16'hd4a4;
assign i[1904]= 16'hd666;
assign i[1905]= 16'hd89e;
assign i[1906]= 16'hdb34;
assign i[1907]= 16'hde13;
assign i[1908]= 16'he122;
assign i[1909]= 16'he44c;
assign i[1910]= 16'he779;
assign i[1911]= 16'hea97;
assign i[1912]= 16'hed91;
assign i[1913]= 16'hf058;
assign i[1914]= 16'hf2dd;
assign i[1915]= 16'hf515;
assign i[1916]= 16'hf6f6;
assign i[1917]= 16'hf87b;
assign i[1918]= 16'hf99e;
assign i[1919]= 16'hfa5d;
assign i[1920]= 16'hfab9;
assign i[1921]= 16'hfab4;
assign i[1922]= 16'hfa53;
assign i[1923]= 16'hf99a;
assign i[1924]= 16'hf892;
assign i[1925]= 16'hf743;
assign i[1926]= 16'hf5b9;
assign i[1927]= 16'hf3ff;
assign i[1928]= 16'hf222;
assign i[1929]= 16'hf031;
assign i[1930]= 16'hee3c;
assign i[1931]= 16'hec52;
assign i[1932]= 16'hea84;
assign i[1933]= 16'he8e3;
assign i[1934]= 16'he780;
assign i[1935]= 16'he66b;
assign i[1936]= 16'he5b5;
assign i[1937]= 16'he56b;
assign i[1938]= 16'he59a;
assign i[1939]= 16'he64c;
assign i[1940]= 16'he788;
assign i[1941]= 16'he953;
assign i[1942]= 16'hebac;
assign i[1943]= 16'hee91;
assign i[1944]= 16'hf1f8;
assign i[1945]= 16'hf5d7;
assign i[1946]= 16'hfa1e;
assign i[1947]= 16'hfeb6;
assign i[1948]= 16'h389;
assign i[1949]= 16'h87e;
assign i[1950]= 16'hd75;
assign i[1951]= 16'h1250;
assign i[1952]= 16'h16ee;
assign i[1953]= 16'h1b31;
assign i[1954]= 16'h1efa;
assign i[1955]= 16'h222c;
assign i[1956]= 16'h24ad;
assign i[1957]= 16'h2669;
assign i[1958]= 16'h274e;
assign i[1959]= 16'h2752;
assign i[1960]= 16'h266e;
assign i[1961]= 16'h24a5;
assign i[1962]= 16'h21fd;
assign i[1963]= 16'h1e83;
assign i[1964]= 16'h1a4a;
assign i[1965]= 16'h156d;
assign i[1966]= 16'h1007;
assign i[1967]= 16'ha3b;
assign i[1968]= 16'h42c;
assign i[1969]= 16'hfe01;
assign i[1970]= 16'hf7e0;
assign i[1971]= 16'hf1f0;
assign i[1972]= 16'hec55;
assign i[1973]= 16'he733;
assign i[1974]= 16'he2a7;
assign i[1975]= 16'hdecd;
assign i[1976]= 16'hdbba;
assign i[1977]= 16'hd97e;
assign i[1978]= 16'hd823;
assign i[1979]= 16'hd7af;
assign i[1980]= 16'hd81f;
assign i[1981]= 16'hd96d;
assign i[1982]= 16'hdb8d;
assign i[1983]= 16'hde6d;
assign i[1984]= 16'he1f9;
assign i[1985]= 16'he619;
assign i[1986]= 16'heab1;
assign i[1987]= 16'hefa5;
assign i[1988]= 16'hf4d6;
assign i[1989]= 16'hfa27;
assign i[1990]= 16'hff7a;
assign i[1991]= 16'h4b0;
assign i[1992]= 16'h9b1;
assign i[1993]= 16'he62;
assign i[1994]= 16'h12ad;
assign i[1995]= 16'h167c;
assign i[1996]= 16'h19bf;
assign i[1997]= 16'h1c67;
assign i[1998]= 16'h1e6a;
assign i[1999]= 16'h1fbe;
assign i[2000]= 16'h2060;
assign i[2001]= 16'h204d;
assign i[2002]= 16'h1f86;
assign i[2003]= 16'h1e11;
assign i[2004]= 16'h1bf4;
assign i[2005]= 16'h1939;
assign i[2006]= 16'h15ed;
assign i[2007]= 16'h1220;
assign i[2008]= 16'hde2;
assign i[2009]= 16'h949;
assign i[2010]= 16'h469;
assign i[2011]= 16'hff5c;
assign i[2012]= 16'hfa3a;
assign i[2013]= 16'hf51c;
assign i[2014]= 16'hf01f;
assign i[2015]= 16'heb5e;
assign i[2016]= 16'he6f3;
assign i[2017]= 16'he2f7;
assign i[2018]= 16'hdf84;
assign i[2019]= 16'hdcae;
assign i[2020]= 16'hda89;
assign i[2021]= 16'hd925;
assign i[2022]= 16'hd88e;
assign i[2023]= 16'hd8ca;
assign i[2024]= 16'hd9dd;
assign i[2025]= 16'hdbc4;
assign i[2026]= 16'hde78;
assign i[2027]= 16'he1ed;
assign i[2028]= 16'he611;
assign i[2029]= 16'head0;
assign i[2030]= 16'hf00f;
assign i[2031]= 16'hf5b3;
assign i[2032]= 16'hfb9b;
assign i[2033]= 16'h1a7;
assign i[2034]= 16'h7b7;
assign i[2035]= 16'hda7;
assign i[2036]= 16'h1359;
assign i[2037]= 16'h18ae;
assign i[2038]= 16'h1d8b;
assign i[2039]= 16'h21d7;
assign i[2040]= 16'h2581;
assign i[2041]= 16'h2879;
assign i[2042]= 16'h2ab5;
assign i[2043]= 16'h2c33;
assign i[2044]= 16'h2cf2;
assign i[2045]= 16'h2cf9;
assign i[2046]= 16'h2c52;
assign i[2047]= 16'h2b0d;
assign i[2048]= 16'h293c;
assign i[2049]= 16'h26f4;
assign i[2050]= 16'h244c;
assign i[2051]= 16'h215e;
assign i[2052]= 16'h1e42;
assign i[2053]= 16'h1b11;
assign i[2054]= 16'h17e3;
assign i[2055]= 16'h14ce;
assign i[2056]= 16'h11e6;
assign i[2057]= 16'hf3b;
assign i[2058]= 16'hcdc;
assign i[2059]= 16'had5;
assign i[2060]= 16'h92b;
assign i[2061]= 16'h7e5;
assign i[2062]= 16'h703;
assign i[2063]= 16'h683;
assign i[2064]= 16'h663;
assign i[2065]= 16'h69b;
assign i[2066]= 16'h723;
assign i[2067]= 16'h7f2;
assign i[2068]= 16'h8fe;
assign i[2069]= 16'ha39;
assign i[2070]= 16'hb9a;
assign i[2071]= 16'hd13;
assign i[2072]= 16'he98;
assign i[2073]= 16'h101d;
assign i[2074]= 16'h1197;
assign i[2075]= 16'h12fa;
assign i[2076]= 16'h143b;
assign i[2077]= 16'h1552;
assign i[2078]= 16'h1634;
assign i[2079]= 16'h16d8;
assign i[2080]= 16'h1739;
assign i[2081]= 16'h174e;
assign i[2082]= 16'h1713;
assign i[2083]= 16'h1684;
assign i[2084]= 16'h159e;
assign i[2085]= 16'h1462;
assign i[2086]= 16'h12d1;
assign i[2087]= 16'h10ee;
assign i[2088]= 16'hec0;
assign i[2089]= 16'hc4f;
assign i[2090]= 16'h9a7;
assign i[2091]= 16'h6d5;
assign i[2092]= 16'h3e8;
assign i[2093]= 16'hf2;
assign i[2094]= 16'hfe08;
assign i[2095]= 16'hfb3d;
assign i[2096]= 16'hf8a6;
assign i[2097]= 16'hf65a;
assign i[2098]= 16'hf46c;
assign i[2099]= 16'hf2f1;
assign i[2100]= 16'hf1f9;
assign i[2101]= 16'hf194;
assign i[2102]= 16'hf1ca;
assign i[2103]= 16'hf2a4;
assign i[2104]= 16'hf423;
assign i[2105]= 16'hf643;
assign i[2106]= 16'hf8fd;
assign i[2107]= 16'hfc42;
assign i[2108]= 16'h0;
assign i[2109]= 16'h41f;
assign i[2110]= 16'h883;
assign i[2111]= 16'hd0e;
assign i[2112]= 16'h119c;
assign i[2113]= 16'h160c;
assign i[2114]= 16'h1a3a;
assign i[2115]= 16'h1e01;
assign i[2116]= 16'h2142;
assign i[2117]= 16'h23de;
assign i[2118]= 16'h25bb;
assign i[2119]= 16'h26c4;
assign i[2120]= 16'h26e9;
assign i[2121]= 16'h2622;
assign i[2122]= 16'h246c;
assign i[2123]= 16'h21cb;
assign i[2124]= 16'h1e4c;
assign i[2125]= 16'h19ff;
assign i[2126]= 16'h14fc;
assign i[2127]= 16'hf5f;
assign i[2128]= 16'h948;
assign i[2129]= 16'h2db;
assign i[2130]= 16'hfc3e;
assign i[2131]= 16'hf593;
assign i[2132]= 16'hef02;
assign i[2133]= 16'he8ad;
assign i[2134]= 16'he2b4;
assign i[2135]= 16'hdd34;
assign i[2136]= 16'hd844;
assign i[2137]= 16'hd3f6;
assign i[2138]= 16'hd056;
assign i[2139]= 16'hcd6b;
assign i[2140]= 16'hcb36;
assign i[2141]= 16'hc9b2;
assign i[2142]= 16'hc8d4;
assign i[2143]= 16'hc88f;
assign i[2144]= 16'hc8d1;
assign i[2145]= 16'hc984;
assign i[2146]= 16'hca90;
assign i[2147]= 16'hcbe0;
assign i[2148]= 16'hcd5a;
assign i[2149]= 16'hcee7;
assign i[2150]= 16'hd073;
assign i[2151]= 16'hd1ea;
assign i[2152]= 16'hd33d;
assign i[2153]= 16'hd460;
assign i[2154]= 16'hd548;
assign i[2155]= 16'hd5f2;
assign i[2156]= 16'hd65b;
assign i[2157]= 16'hd687;
assign i[2158]= 16'hd67a;
assign i[2159]= 16'hd63b;
assign i[2160]= 16'hd5d5;
assign i[2161]= 16'hd554;
assign i[2162]= 16'hd4c4;
assign i[2163]= 16'hd432;
assign i[2164]= 16'hd3ab;
assign i[2165]= 16'hd33b;
assign i[2166]= 16'hd2ee;
assign i[2167]= 16'hd2cc;
assign i[2168]= 16'hd2df;
assign i[2169]= 16'hd32c;
assign i[2170]= 16'hd3b8;
assign i[2171]= 16'hd484;
assign i[2172]= 16'hd592;
assign i[2173]= 16'hd6e0;
assign i[2174]= 16'hd86b;
assign i[2175]= 16'hda30;
assign i[2176]= 16'hdc28;
assign i[2177]= 16'hde50;
assign i[2178]= 16'he09f;
assign i[2179]= 16'he310;
assign i[2180]= 16'he59b;
assign i[2181]= 16'he83b;
assign i[2182]= 16'heae9;
assign i[2183]= 16'hed9e;
assign i[2184]= 16'hf054;
assign i[2185]= 16'hf306;
assign i[2186]= 16'hf5ad;
assign i[2187]= 16'hf845;
assign i[2188]= 16'hfac9;
assign i[2189]= 16'hfd32;
assign i[2190]= 16'hff7d;
assign i[2191]= 16'h1a3;
assign i[2192]= 16'h3a1;
assign i[2193]= 16'h572;
assign i[2194]= 16'h710;
assign i[2195]= 16'h878;
assign i[2196]= 16'h9a5;
assign i[2197]= 16'ha94;
assign i[2198]= 16'hb41;
assign i[2199]= 16'hbaa;
assign i[2200]= 16'hbce;
assign i[2201]= 16'hbac;
assign i[2202]= 16'hb45;
assign i[2203]= 16'ha9a;
assign i[2204]= 16'h9ad;
assign i[2205]= 16'h883;
assign i[2206]= 16'h721;
assign i[2207]= 16'h58c;
assign i[2208]= 16'h3cc;
assign i[2209]= 16'h1e7;
assign i[2210]= 16'hffe8;
assign i[2211]= 16'hfdd5;
assign i[2212]= 16'hfbb8;
assign i[2213]= 16'hf999;
assign i[2214]= 16'hf782;
assign i[2215]= 16'hf57c;
assign i[2216]= 16'hf38e;
assign i[2217]= 16'hf1c0;
assign i[2218]= 16'hf019;
assign i[2219]= 16'heea0;
assign i[2220]= 16'hed5a;
assign i[2221]= 16'hec4b;
assign i[2222]= 16'heb79;
assign i[2223]= 16'heae5;
assign i[2224]= 16'hea92;
assign i[2225]= 16'hea82;
assign i[2226]= 16'heab4;
assign i[2227]= 16'heb2a;
assign i[2228]= 16'hebe2;
assign i[2229]= 16'hecd9;
assign i[2230]= 16'hee0e;
assign i[2231]= 16'hef7d;
assign i[2232]= 16'hf120;
assign i[2233]= 16'hf2f3;
assign i[2234]= 16'hf4f0;
assign i[2235]= 16'hf70d;
assign i[2236]= 16'hf945;
assign i[2237]= 16'hfb8c;
assign i[2238]= 16'hfddb;
assign i[2239]= 16'h25;
assign i[2240]= 16'h262;
assign i[2241]= 16'h487;
assign i[2242]= 16'h689;
assign i[2243]= 16'h860;
assign i[2244]= 16'ha02;
assign i[2245]= 16'hb68;
assign i[2246]= 16'hc8e;
assign i[2247]= 16'hd6e;
assign i[2248]= 16'he09;
assign i[2249]= 16'he5f;
assign i[2250]= 16'he73;
assign i[2251]= 16'he4d;
assign i[2252]= 16'hdf6;
assign i[2253]= 16'hd78;
assign i[2254]= 16'hce0;
assign i[2255]= 16'hc3f;
assign i[2256]= 16'hba4;
assign i[2257]= 16'hb21;
assign i[2258]= 16'hac5;
assign i[2259]= 16'haa1;
assign i[2260]= 16'hac3;
assign i[2261]= 16'hb37;
assign i[2262]= 16'hc08;
assign i[2263]= 16'hd3a;
assign i[2264]= 16'hecf;
assign i[2265]= 16'h10c5;
assign i[2266]= 16'h1314;
assign i[2267]= 16'h15b2;
assign i[2268]= 16'h188d;
assign i[2269]= 16'h1b92;
assign i[2270]= 16'h1ea9;
assign i[2271]= 16'h21b8;
assign i[2272]= 16'h24a1;
assign i[2273]= 16'h2747;
assign i[2274]= 16'h298c;
assign i[2275]= 16'h2b54;
assign i[2276]= 16'h2c85;
assign i[2277]= 16'h2d08;
assign i[2278]= 16'h2cca;
assign i[2279]= 16'h2bbe;
assign i[2280]= 16'h29dd;
assign i[2281]= 16'h2725;
assign i[2282]= 16'h239c;
assign i[2283]= 16'h1f50;
assign i[2284]= 16'h1a53;
assign i[2285]= 16'h14be;
assign i[2286]= 16'heb1;
assign i[2287]= 16'h84f;
assign i[2288]= 16'h1be;
assign i[2289]= 16'hfb29;
assign i[2290]= 16'hf4b7;
assign i[2291]= 16'hee94;
assign i[2292]= 16'he8e7;
assign i[2293]= 16'he3d5;
assign i[2294]= 16'hdf7f;
assign i[2295]= 16'hdbfe;
assign i[2296]= 16'hd967;
assign i[2297]= 16'hd7c9;
assign i[2298]= 16'hd729;
assign i[2299]= 16'hd787;
assign i[2300]= 16'hd8d8;
assign i[2301]= 16'hdb0e;
assign i[2302]= 16'hde13;
assign i[2303]= 16'he1cc;
assign i[2304]= 16'he617;
assign i[2305]= 16'head4;
assign i[2306]= 16'hefdb;
assign i[2307]= 16'hf509;
assign i[2308]= 16'hfa36;
assign i[2309]= 16'hff42;
assign i[2310]= 16'h409;
assign i[2311]= 16'h872;
assign i[2312]= 16'hc65;
assign i[2313]= 16'hfcf;
assign i[2314]= 16'h12a4;
assign i[2315]= 16'h14dd;
assign i[2316]= 16'h167a;
assign i[2317]= 16'h177e;
assign i[2318]= 16'h17f4;
assign i[2319]= 16'h17e7;
assign i[2320]= 16'h1769;
assign i[2321]= 16'h168d;
assign i[2322]= 16'h1565;
assign i[2323]= 16'h1407;
assign i[2324]= 16'h1285;
assign i[2325]= 16'h10f3;
assign i[2326]= 16'hf5f;
assign i[2327]= 16'hdd5;
assign i[2328]= 16'hc60;
assign i[2329]= 16'hb05;
assign i[2330]= 16'h9c6;
assign i[2331]= 16'h8a1;
assign i[2332]= 16'h791;
assign i[2333]= 16'h68f;
assign i[2334]= 16'h590;
assign i[2335]= 16'h48a;
assign i[2336]= 16'h36f;
assign i[2337]= 16'h234;
assign i[2338]= 16'hcd;
assign i[2339]= 16'hff32;
assign i[2340]= 16'hfd57;
assign i[2341]= 16'hfb3b;
assign i[2342]= 16'hf8da;
assign i[2343]= 16'hf636;
assign i[2344]= 16'hf354;
assign i[2345]= 16'hf03f;
assign i[2346]= 16'hed00;
assign i[2347]= 16'he9a8;
assign i[2348]= 16'he649;
assign i[2349]= 16'he2f7;
assign i[2350]= 16'hdfc6;
assign i[2351]= 16'hdccc;
assign i[2352]= 16'hda20;
assign i[2353]= 16'hd7d7;
assign i[2354]= 16'hd603;
assign i[2355]= 16'hd4b6;
assign i[2356]= 16'hd3ff;
assign i[2357]= 16'hd3e9;
assign i[2358]= 16'hd47c;
assign i[2359]= 16'hd5bd;
assign i[2360]= 16'hd7aa;
assign i[2361]= 16'hda40;
assign i[2362]= 16'hdd78;
assign i[2363]= 16'he147;
assign i[2364]= 16'he59e;
assign i[2365]= 16'hea6b;
assign i[2366]= 16'hef9b;
assign i[2367]= 16'hf518;
assign i[2368]= 16'hfacb;
assign i[2369]= 16'h9c;
assign i[2370]= 16'h672;
assign i[2371]= 16'hc36;
assign i[2372]= 16'h11d0;
assign i[2373]= 16'h1728;
assign i[2374]= 16'h1c29;
assign i[2375]= 16'h20bf;
assign i[2376]= 16'h24d9;
assign i[2377]= 16'h2866;
assign i[2378]= 16'h2b5a;
assign i[2379]= 16'h2da9;
assign i[2380]= 16'h2f4c;
assign i[2381]= 16'h303c;
assign i[2382]= 16'h3076;
assign i[2383]= 16'h2ffa;
assign i[2384]= 16'h2ecb;
assign i[2385]= 16'h2cee;
assign i[2386]= 16'h2a6a;
assign i[2387]= 16'h2749;
assign i[2388]= 16'h2399;
assign i[2389]= 16'h1f67;
assign i[2390]= 16'h1ac5;
assign i[2391]= 16'h15c5;
assign i[2392]= 16'h107c;
assign i[2393]= 16'hb00;
assign i[2394]= 16'h567;
assign i[2395]= 16'hffcb;
assign i[2396]= 16'hfa40;
assign i[2397]= 16'hf4df;
assign i[2398]= 16'hefbf;
assign i[2399]= 16'heaf7;
assign i[2400]= 16'he699;
assign i[2401]= 16'he2ba;
assign i[2402]= 16'hdf68;
assign i[2403]= 16'hdcb0;
assign i[2404]= 16'hda9e;
assign i[2405]= 16'hd937;
assign i[2406]= 16'hd87f;
assign i[2407]= 16'hd874;
assign i[2408]= 16'hd914;
assign i[2409]= 16'hda55;
assign i[2410]= 16'hdc2c;
assign i[2411]= 16'hde8c;
assign i[2412]= 16'he161;
assign i[2413]= 16'he499;
assign i[2414]= 16'he81c;
assign i[2415]= 16'hebd5;
assign i[2416]= 16'hefa9;
assign i[2417]= 16'hf380;
assign i[2418]= 16'hf742;
assign i[2419]= 16'hfad5;
assign i[2420]= 16'hfe24;
assign i[2421]= 16'h118;
assign i[2422]= 16'h3a0;
assign i[2423]= 16'h5ab;
assign i[2424]= 16'h72b;
assign i[2425]= 16'h816;
assign i[2426]= 16'h864;
assign i[2427]= 16'h811;
assign i[2428]= 16'h71d;
assign i[2429]= 16'h58a;
assign i[2430]= 16'h35e;
assign i[2431]= 16'ha2;
assign i[2432]= 16'hfd62;
assign i[2433]= 16'hf9a9;
assign i[2434]= 16'hf58a;
assign i[2435]= 16'hf117;
assign i[2436]= 16'hec64;
assign i[2437]= 16'he785;
assign i[2438]= 16'he292;
assign i[2439]= 16'hdda2;
assign i[2440]= 16'hd8cc;
assign i[2441]= 16'hd428;
assign i[2442]= 16'hcfcd;
assign i[2443]= 16'hcbd2;
assign i[2444]= 16'hc84b;
assign i[2445]= 16'hc54e;
assign i[2446]= 16'hc2ed;
assign i[2447]= 16'hc136;
assign i[2448]= 16'hc03a;
assign i[2449]= 16'hc002;
assign i[2450]= 16'hc093;
assign i[2451]= 16'hc1f4;
assign i[2452]= 16'hc426;
assign i[2453]= 16'hc722;
assign i[2454]= 16'hcae2;
assign i[2455]= 16'hcf5a;
assign i[2456]= 16'hd479;
assign i[2457]= 16'hda2b;
assign i[2458]= 16'he057;
assign i[2459]= 16'he6e3;
assign i[2460]= 16'hedaf;
assign i[2461]= 16'hf49c;
assign i[2462]= 16'hfb86;
assign i[2463]= 16'h248;
assign i[2464]= 16'h8c2;
assign i[2465]= 16'hed0;
assign i[2466]= 16'h144f;
assign i[2467]= 16'h1922;
assign i[2468]= 16'h1d2d;
assign i[2469]= 16'h205a;
assign i[2470]= 16'h2295;
assign i[2471]= 16'h23d2;
assign i[2472]= 16'h240c;
assign i[2473]= 16'h2340;
assign i[2474]= 16'h2177;
assign i[2475]= 16'h1ebb;
assign i[2476]= 16'h1b20;
assign i[2477]= 16'h16bf;
assign i[2478]= 16'h11b4;
assign i[2479]= 16'hc23;
assign i[2480]= 16'h62f;
assign i[2481]= 16'h2;
assign i[2482]= 16'hf9c6;
assign i[2483]= 16'hf3a3;
assign i[2484]= 16'hedc1;
assign i[2485]= 16'he848;
assign i[2486]= 16'he35b;
assign i[2487]= 16'hdf1b;
assign i[2488]= 16'hdba1;
assign i[2489]= 16'hd903;
assign i[2490]= 16'hd750;
assign i[2491]= 16'hd690;
assign i[2492]= 16'hd6c7;
assign i[2493]= 16'hd7f0;
assign i[2494]= 16'hda00;
assign i[2495]= 16'hdce9;
assign i[2496]= 16'he096;
assign i[2497]= 16'he4ec;
assign i[2498]= 16'he9d1;
assign i[2499]= 16'hef26;
assign i[2500]= 16'hf4ca;
assign i[2501]= 16'hfa9c;
assign i[2502]= 16'h7c;
assign i[2503]= 16'h64d;
assign i[2504]= 16'hbf1;
assign i[2505]= 16'h114f;
assign i[2506]= 16'h1650;
assign i[2507]= 16'h1ae3;
assign i[2508]= 16'h1ef8;
assign i[2509]= 16'h2285;
assign i[2510]= 16'h2585;
assign i[2511]= 16'h27f6;
assign i[2512]= 16'h29d9;
assign i[2513]= 16'h2b34;
assign i[2514]= 16'h2c0d;
assign i[2515]= 16'h2c6f;
assign i[2516]= 16'h2c65;
assign i[2517]= 16'h2bfd;
assign i[2518]= 16'h2b43;
assign i[2519]= 16'h2a45;
assign i[2520]= 16'h2911;
assign i[2521]= 16'h27b2;
assign i[2522]= 16'h2634;
assign i[2523]= 16'h24a2;
assign i[2524]= 16'h2305;
assign i[2525]= 16'h2165;
assign i[2526]= 16'h1fc8;
assign i[2527]= 16'h1e34;
assign i[2528]= 16'h1cae;
assign i[2529]= 16'h1b3a;
assign i[2530]= 16'h19dc;
assign i[2531]= 16'h1897;
assign i[2532]= 16'h176e;
assign i[2533]= 16'h1665;
assign i[2534]= 16'h1580;
assign i[2535]= 16'h14c2;
assign i[2536]= 16'h142f;
assign i[2537]= 16'h13cd;
assign i[2538]= 16'h139f;
assign i[2539]= 16'h13ab;
assign i[2540]= 16'h13f3;
assign i[2541]= 16'h147c;
assign i[2542]= 16'h1548;
assign i[2543]= 16'h165a;
assign i[2544]= 16'h17b0;
assign i[2545]= 16'h194a;
assign i[2546]= 16'h1b26;
assign i[2547]= 16'h1d3c;
assign i[2548]= 16'h1f87;
assign i[2549]= 16'h21fe;
assign i[2550]= 16'h2495;
assign i[2551]= 16'h2740;
assign i[2552]= 16'h29f1;
assign i[2553]= 16'h2c98;
assign i[2554]= 16'h2f24;
assign i[2555]= 16'h3185;
assign i[2556]= 16'h33ab;
assign i[2557]= 16'h3584;
assign i[2558]= 16'h3701;
assign i[2559]= 16'h3814;
assign i[2560]= 16'h38b1;
assign i[2561]= 16'h38cd;
assign i[2562]= 16'h3861;
assign i[2563]= 16'h3766;
assign i[2564]= 16'h35da;
assign i[2565]= 16'h33bd;
assign i[2566]= 16'h3113;
assign i[2567]= 16'h2de1;
assign i[2568]= 16'h2a2f;
assign i[2569]= 16'h2608;
assign i[2570]= 16'h2179;
assign i[2571]= 16'h1c91;
assign i[2572]= 16'h175f;
assign i[2573]= 16'h11f4;
assign i[2574]= 16'hc63;
assign i[2575]= 16'h6bd;
assign i[2576]= 16'h115;
assign i[2577]= 16'hfb7e;
assign i[2578]= 16'hf607;
assign i[2579]= 16'hf0c1;
assign i[2580]= 16'hebbe;
assign i[2581]= 16'he70a;
assign i[2582]= 16'he2b5;
assign i[2583]= 16'hdec9;
assign i[2584]= 16'hdb52;
assign i[2585]= 16'hd85a;
assign i[2586]= 16'hd5e8;
assign i[2587]= 16'hd403;
assign i[2588]= 16'hd2b2;
assign i[2589]= 16'hd1f6;
assign i[2590]= 16'hd1d4;
assign i[2591]= 16'hd24b;
assign i[2592]= 16'hd35c;
assign i[2593]= 16'hd504;
assign i[2594]= 16'hd73f;
assign i[2595]= 16'hda07;
assign i[2596]= 16'hdd53;
assign i[2597]= 16'he11c;
assign i[2598]= 16'he554;
assign i[2599]= 16'he9ed;
assign i[2600]= 16'heed9;
assign i[2601]= 16'hf405;
assign i[2602]= 16'hf95d;
assign i[2603]= 16'hfece;
assign i[2604]= 16'h441;
assign i[2605]= 16'h99f;
assign i[2606]= 16'hed1;
assign i[2607]= 16'h13c1;
assign i[2608]= 16'h1856;
assign i[2609]= 16'h1c7d;
assign i[2610]= 16'h2020;
assign i[2611]= 16'h232f;
assign i[2612]= 16'h259b;
assign i[2613]= 16'h2759;
assign i[2614]= 16'h2860;
assign i[2615]= 16'h28ad;
assign i[2616]= 16'h2841;
assign i[2617]= 16'h2720;
assign i[2618]= 16'h2554;
assign i[2619]= 16'h22eb;
assign i[2620]= 16'h1ff5;
assign i[2621]= 16'h1c88;
assign i[2622]= 16'h18bc;
assign i[2623]= 16'h14ab;
assign i[2624]= 16'h1072;
assign i[2625]= 16'hc2d;
assign i[2626]= 16'h7fa;
assign i[2627]= 16'h3f4;
assign i[2628]= 16'h37;
assign i[2629]= 16'hfcda;
assign i[2630]= 16'hf9f2;
assign i[2631]= 16'hf78f;
assign i[2632]= 16'hf5bf;
assign i[2633]= 16'hf489;
assign i[2634]= 16'hf3ef;
assign i[2635]= 16'hf3f1;
assign i[2636]= 16'hf486;
assign i[2637]= 16'hf5a3;
assign i[2638]= 16'hf738;
assign i[2639]= 16'hf930;
assign i[2640]= 16'hfb75;
assign i[2641]= 16'hfdef;
assign i[2642]= 16'h81;
assign i[2643]= 16'h314;
assign i[2644]= 16'h58d;
assign i[2645]= 16'h7d2;
assign i[2646]= 16'h9ce;
assign i[2647]= 16'hb6d;
assign i[2648]= 16'hca0;
assign i[2649]= 16'hd5c;
assign i[2650]= 16'hd99;
assign i[2651]= 16'hd55;
assign i[2652]= 16'hc92;
assign i[2653]= 16'hb58;
assign i[2654]= 16'h9b1;
assign i[2655]= 16'h7ac;
assign i[2656]= 16'h559;
assign i[2657]= 16'h2ce;
assign i[2658]= 16'h20;
assign i[2659]= 16'hfd64;
assign i[2660]= 16'hfab0;
assign i[2661]= 16'hf818;
assign i[2662]= 16'hf5ae;
assign i[2663]= 16'hf384;
assign i[2664]= 16'hf1a6;
assign i[2665]= 16'hf01d;
assign i[2666]= 16'heeef;
assign i[2667]= 16'hee1d;
assign i[2668]= 16'heda6;
assign i[2669]= 16'hed82;
assign i[2670]= 16'heda8;
assign i[2671]= 16'hee0d;
assign i[2672]= 16'heea1;
assign i[2673]= 16'hef54;
assign i[2674]= 16'hf015;
assign i[2675]= 16'hf0d5;
assign i[2676]= 16'hf183;
assign i[2677]= 16'hf210;
assign i[2678]= 16'hf272;
assign i[2679]= 16'hf2a0;
assign i[2680]= 16'hf293;
assign i[2681]= 16'hf24b;
assign i[2682]= 16'hf1ca;
assign i[2683]= 16'hf115;
assign i[2684]= 16'hf037;
assign i[2685]= 16'hef3c;
assign i[2686]= 16'hee36;
assign i[2687]= 16'hed35;
assign i[2688]= 16'hec4e;
assign i[2689]= 16'heb95;
assign i[2690]= 16'heb1d;
assign i[2691]= 16'heafb;
assign i[2692]= 16'heb3f;
assign i[2693]= 16'hebf7;
assign i[2694]= 16'hed2d;
assign i[2695]= 16'heee9;
assign i[2696]= 16'hf12d;
assign i[2697]= 16'hf3f6;
assign i[2698]= 16'hf73c;
assign i[2699]= 16'hfaf3;
assign i[2700]= 16'hff0a;
assign i[2701]= 16'h36c;
assign i[2702]= 16'h800;
assign i[2703]= 16'hcac;
assign i[2704]= 16'h1152;
assign i[2705]= 16'h15d4;
assign i[2706]= 16'h1a14;
assign i[2707]= 16'h1df4;
assign i[2708]= 16'h215b;
assign i[2709]= 16'h2430;
assign i[2710]= 16'h265f;
assign i[2711]= 16'h27d8;
assign i[2712]= 16'h2890;
assign i[2713]= 16'h2884;
assign i[2714]= 16'h27b2;
assign i[2715]= 16'h2622;
assign i[2716]= 16'h23de;
assign i[2717]= 16'h20f7;
assign i[2718]= 16'h1d81;
assign i[2719]= 16'h1996;
assign i[2720]= 16'h1551;
assign i[2721]= 16'h10cf;
assign i[2722]= 16'hc2f;
assign i[2723]= 16'h78f;
assign i[2724]= 16'h30b;
assign i[2725]= 16'hfec1;
assign i[2726]= 16'hfac5;
assign i[2727]= 16'hf72f;
assign i[2728]= 16'hf40d;
assign i[2729]= 16'hf16c;
assign i[2730]= 16'hef51;
assign i[2731]= 16'hedbe;
assign i[2732]= 16'hecaf;
assign i[2733]= 16'hec1c;
assign i[2734]= 16'hebf7;
assign i[2735]= 16'hec31;
assign i[2736]= 16'hecb6;
assign i[2737]= 16'hed70;
assign i[2738]= 16'hee49;
assign i[2739]= 16'hef2a;
assign i[2740]= 16'heffc;
assign i[2741]= 16'hf0ab;
assign i[2742]= 16'hf123;
assign i[2743]= 16'hf155;
assign i[2744]= 16'hf135;
assign i[2745]= 16'hf0bb;
assign i[2746]= 16'hefe2;
assign i[2747]= 16'heeab;
assign i[2748]= 16'hed1a;
assign i[2749]= 16'heb38;
assign i[2750]= 16'he910;
assign i[2751]= 16'he6b0;
assign i[2752]= 16'he42a;
assign i[2753]= 16'he18f;
assign i[2754]= 16'hdef4;
assign i[2755]= 16'hdc69;
assign i[2756]= 16'hda02;
assign i[2757]= 16'hd7ce;
assign i[2758]= 16'hd5da;
assign i[2759]= 16'hd433;
assign i[2760]= 16'hd2df;
assign i[2761]= 16'hd1e2;
assign i[2762]= 16'hd13c;
assign i[2763]= 16'hd0e9;
assign i[2764]= 16'hd0e2;
assign i[2765]= 16'hd11d;
assign i[2766]= 16'hd18c;
assign i[2767]= 16'hd221;
assign i[2768]= 16'hd2cc;
assign i[2769]= 16'hd37c;
assign i[2770]= 16'hd41f;
assign i[2771]= 16'hd4a8;
assign i[2772]= 16'hd507;
assign i[2773]= 16'hd533;
assign i[2774]= 16'hd523;
assign i[2775]= 16'hd4d3;
assign i[2776]= 16'hd442;
assign i[2777]= 16'hd375;
assign i[2778]= 16'hd272;
assign i[2779]= 16'hd145;
assign i[2780]= 16'hcffd;
assign i[2781]= 16'hceac;
assign i[2782]= 16'hcd67;
assign i[2783]= 16'hcc43;
assign i[2784]= 16'hcb56;
assign i[2785]= 16'hcab8;
assign i[2786]= 16'hca7e;
assign i[2787]= 16'hcabb;
assign i[2788]= 16'hcb81;
assign i[2789]= 16'hccdd;
assign i[2790]= 16'hced8;
assign i[2791]= 16'hd177;
assign i[2792]= 16'hd4bb;
assign i[2793]= 16'hd89e;
assign i[2794]= 16'hdd17;
assign i[2795]= 16'he216;
assign i[2796]= 16'he78a;
assign i[2797]= 16'hed5a;
assign i[2798]= 16'hf36c;
assign i[2799]= 16'hf9a4;
assign i[2800]= 16'hffe3;
assign i[2801]= 16'h60a;
assign i[2802]= 16'hbf9;
assign i[2803]= 16'h1194;
assign i[2804]= 16'h16bd;
assign i[2805]= 16'h1b5b;
assign i[2806]= 16'h1f56;
assign i[2807]= 16'h229d;
assign i[2808]= 16'h2521;
assign i[2809]= 16'h26d8;
assign i[2810]= 16'h27bd;
assign i[2811]= 16'h27cf;
assign i[2812]= 16'h2711;
assign i[2813]= 16'h258c;
assign i[2814]= 16'h234a;
assign i[2815]= 16'h205c;
assign i[2816]= 16'h1cd2;
assign i[2817]= 16'h18c1;
assign i[2818]= 16'h143f;
assign i[2819]= 16'hf62;
assign i[2820]= 16'ha41;
assign i[2821]= 16'h4f5;
assign i[2822]= 16'hff94;
assign i[2823]= 16'hfa33;
assign i[2824]= 16'hf4e8;
assign i[2825]= 16'hefc6;
assign i[2826]= 16'heae0;
assign i[2827]= 16'he645;
assign i[2828]= 16'he205;
assign i[2829]= 16'hde2c;
assign i[2830]= 16'hdac5;
assign i[2831]= 16'hd7da;
assign i[2832]= 16'hd572;
assign i[2833]= 16'hd393;
assign i[2834]= 16'hd242;
assign i[2835]= 16'hd181;
assign i[2836]= 16'hd151;
assign i[2837]= 16'hd1b1;
assign i[2838]= 16'hd29d;
assign i[2839]= 16'hd413;
assign i[2840]= 16'hd60a;
assign i[2841]= 16'hd87b;
assign i[2842]= 16'hdb59;
assign i[2843]= 16'hde9a;
assign i[2844]= 16'he22c;
assign i[2845]= 16'he600;
assign i[2846]= 16'hea04;
assign i[2847]= 16'hee22;
assign i[2848]= 16'hf247;
assign i[2849]= 16'hf65c;
assign i[2850]= 16'hfa4d;
assign i[2851]= 16'hfe02;
assign i[2852]= 16'h169;
assign i[2853]= 16'h46e;
assign i[2854]= 16'h702;
assign i[2855]= 16'h916;
assign i[2856]= 16'haa1;
assign i[2857]= 16'hb9b;
assign i[2858]= 16'hc03;
assign i[2859]= 16'hbda;
assign i[2860]= 16'hb26;
assign i[2861]= 16'h9f1;
assign i[2862]= 16'h84a;
assign i[2863]= 16'h643;
assign i[2864]= 16'h3ef;
assign i[2865]= 16'h166;
assign i[2866]= 16'hfec0;
assign i[2867]= 16'hfc14;
assign i[2868]= 16'hf97c;
assign i[2869]= 16'hf70d;
assign i[2870]= 16'hf4dc;
assign i[2871]= 16'hf2fa;
assign i[2872]= 16'hf174;
assign i[2873]= 16'hf052;
assign i[2874]= 16'hef99;
assign i[2875]= 16'hef46;
assign i[2876]= 16'hef54;
assign i[2877]= 16'hefb5;
assign i[2878]= 16'hf05c;
assign i[2879]= 16'hf133;
assign i[2880]= 16'hf225;
assign i[2881]= 16'hf319;
assign i[2882]= 16'hf3f5;
assign i[2883]= 16'hf4a2;
assign i[2884]= 16'hf507;
assign i[2885]= 16'hf510;
assign i[2886]= 16'hf4ac;
assign i[2887]= 16'hf3d0;
assign i[2888]= 16'hf276;
assign i[2889]= 16'hf09d;
assign i[2890]= 16'hee4b;
assign i[2891]= 16'heb8e;
assign i[2892]= 16'he878;
assign i[2893]= 16'he522;
assign i[2894]= 16'he1aa;
assign i[2895]= 16'hde31;
assign i[2896]= 16'hdadb;
assign i[2897]= 16'hd7cd;
assign i[2898]= 16'hd52d;
assign i[2899]= 16'hd31d;
assign i[2900]= 16'hd1bf;
assign i[2901]= 16'hd12d;
assign i[2902]= 16'hd17e;
assign i[2903]= 16'hd2be;
assign i[2904]= 16'hd4f6;
assign i[2905]= 16'hd823;
assign i[2906]= 16'hdc3a;
assign i[2907]= 16'he129;
assign i[2908]= 16'he6d5;
assign i[2909]= 16'hed1b;
assign i[2910]= 16'hf3d2;
assign i[2911]= 16'hfacc;
assign i[2912]= 16'h1d6;
assign i[2913]= 16'h8c0;
assign i[2914]= 16'hf55;
assign i[2915]= 16'h1563;
assign i[2916]= 16'h1abc;
assign i[2917]= 16'h1f37;
assign i[2918]= 16'h22b0;
assign i[2919]= 16'h250e;
assign i[2920]= 16'h263e;
assign i[2921]= 16'h2637;
assign i[2922]= 16'h24fa;
assign i[2923]= 16'h2290;
assign i[2924]= 16'h1f0e;
assign i[2925]= 16'h1a90;
assign i[2926]= 16'h1538;
assign i[2927]= 16'hf30;
assign i[2928]= 16'h8a6;
assign i[2929]= 16'h1cc;
assign i[2930]= 16'hfad5;
assign i[2931]= 16'hf3f0;
assign i[2932]= 16'hed4f;
assign i[2933]= 16'he71e;
assign i[2934]= 16'he183;
assign i[2935]= 16'hdca0;
assign i[2936]= 16'hd88f;
assign i[2937]= 16'hd561;
assign i[2938]= 16'hd31f;
assign i[2939]= 16'hd1cc;
assign i[2940]= 16'hd162;
assign i[2941]= 16'hd1d2;
assign i[2942]= 16'hd308;
assign i[2943]= 16'hd4eb;
assign i[2944]= 16'hd75e;
assign i[2945]= 16'hda40;
assign i[2946]= 16'hdd6e;
assign i[2947]= 16'he0c6;
assign i[2948]= 16'he427;
assign i[2949]= 16'he772;
assign i[2950]= 16'hea8c;
assign i[2951]= 16'hed5c;
assign i[2952]= 16'hefd0;
assign i[2953]= 16'hf1dc;
assign i[2954]= 16'hf378;
assign i[2955]= 16'hf4a2;
assign i[2956]= 16'hf55c;
assign i[2957]= 16'hf5af;
assign i[2958]= 16'hf5a7;
assign i[2959]= 16'hf553;
assign i[2960]= 16'hf4c6;
assign i[2961]= 16'hf413;
assign i[2962]= 16'hf34f;
assign i[2963]= 16'hf28d;
assign i[2964]= 16'hf1e0;
assign i[2965]= 16'hf15b;
assign i[2966]= 16'hf10b;
assign i[2967]= 16'hf0fc;
assign i[2968]= 16'hf138;
assign i[2969]= 16'hf1c2;
assign i[2970]= 16'hf29d;
assign i[2971]= 16'hf3c6;
assign i[2972]= 16'hf538;
assign i[2973]= 16'hf6eb;
assign i[2974]= 16'hf8d6;
assign i[2975]= 16'hfaea;
assign i[2976]= 16'hfd1c;
assign i[2977]= 16'hff5b;
assign i[2978]= 16'h199;
assign i[2979]= 16'h3c9;
assign i[2980]= 16'h5db;
assign i[2981]= 16'h7c3;
assign i[2982]= 16'h974;
assign i[2983]= 16'hae5;
assign i[2984]= 16'hc0c;
assign i[2985]= 16'hce3;
assign i[2986]= 16'hd65;
assign i[2987]= 16'hd8d;
assign i[2988]= 16'hd5a;
assign i[2989]= 16'hccb;
assign i[2990]= 16'hbe1;
assign i[2991]= 16'ha9d;
assign i[2992]= 16'h903;
assign i[2993]= 16'h716;
assign i[2994]= 16'h4db;
assign i[2995]= 16'h257;
assign i[2996]= 16'hff93;
assign i[2997]= 16'hfc93;
assign i[2998]= 16'hf961;
assign i[2999]= 16'hf606;
assign i[3000]= 16'hf28d;
assign i[3001]= 16'hef01;
assign i[3002]= 16'heb6e;
assign i[3003]= 16'he7e3;
assign i[3004]= 16'he46d;
assign i[3005]= 16'he11c;
assign i[3006]= 16'hde00;
assign i[3007]= 16'hdb29;
assign i[3008]= 16'hd8a8;
assign i[3009]= 16'hd68d;
assign i[3010]= 16'hd4e8;
assign i[3011]= 16'hd3c6;
assign i[3012]= 16'hd333;
assign i[3013]= 16'hd33b;
assign i[3014]= 16'hd3e6;
assign i[3015]= 16'hd537;
assign i[3016]= 16'hd732;
assign i[3017]= 16'hd9d4;
assign i[3018]= 16'hdd18;
assign i[3019]= 16'he0f5;
assign i[3020]= 16'he55f;
assign i[3021]= 16'hea47;
assign i[3022]= 16'hef99;
assign i[3023]= 16'hf540;
assign i[3024]= 16'hfb26;
assign i[3025]= 16'h12f;
assign i[3026]= 16'h745;
assign i[3027]= 16'hd4c;
assign i[3028]= 16'h132c;
assign i[3029]= 16'h18cd;
assign i[3030]= 16'h1e18;
assign i[3031]= 16'h22fa;
assign i[3032]= 16'h2763;
assign i[3033]= 16'h2b46;
assign i[3034]= 16'h2e99;
assign i[3035]= 16'h3156;
assign i[3036]= 16'h337d;
assign i[3037]= 16'h350e;
assign i[3038]= 16'h360f;
assign i[3039]= 16'h368a;
assign i[3040]= 16'h3688;
assign i[3041]= 16'h3617;
assign i[3042]= 16'h3547;
assign i[3043]= 16'h3427;
assign i[3044]= 16'h32c7;
assign i[3045]= 16'h3137;
assign i[3046]= 16'h2f85;
assign i[3047]= 16'h2dc1;
assign i[3048]= 16'h2bf4;
assign i[3049]= 16'h2a2a;
assign i[3050]= 16'h2868;
assign i[3051]= 16'h26b5;
assign i[3052]= 16'h2512;
assign i[3053]= 16'h2380;
assign i[3054]= 16'h21fb;
assign i[3055]= 16'h2082;
assign i[3056]= 16'h1f0d;
assign i[3057]= 16'h1d98;
assign i[3058]= 16'h1c1a;
assign i[3059]= 16'h1a8e;
assign i[3060]= 16'h18ec;
assign i[3061]= 16'h172f;
assign i[3062]= 16'h1553;
assign i[3063]= 16'h1355;
assign i[3064]= 16'h1134;
assign i[3065]= 16'hef2;
assign i[3066]= 16'hc91;
assign i[3067]= 16'ha17;
assign i[3068]= 16'h78b;
assign i[3069]= 16'h4f6;
assign i[3070]= 16'h263;
assign i[3071]= 16'hffde;
assign i[3072]= 16'hfd71;
assign i[3073]= 16'hfb2a;
assign i[3074]= 16'hf916;
assign i[3075]= 16'hf740;
assign i[3076]= 16'hf5b3;
assign i[3077]= 16'hf478;
assign i[3078]= 16'hf397;
assign i[3079]= 16'hf314;
assign i[3080]= 16'hf2f2;
assign i[3081]= 16'hf333;
assign i[3082]= 16'hf3d2;
assign i[3083]= 16'hf4cd;
assign i[3084]= 16'hf61b;
assign i[3085]= 16'hf7b3;
assign i[3086]= 16'hf98a;
assign i[3087]= 16'hfb94;
assign i[3088]= 16'hfdc1;
assign i[3089]= 16'h3;
assign i[3090]= 16'h24c;
assign i[3091]= 16'h48d;
assign i[3092]= 16'h6b8;
assign i[3093]= 16'h8bf;
assign i[3094]= 16'ha98;
assign i[3095]= 16'hc3a;
assign i[3096]= 16'hd9c;
assign i[3097]= 16'hebc;
assign i[3098]= 16'hf96;
assign i[3099]= 16'h102b;
assign i[3100]= 16'h1080;
assign i[3101]= 16'h109a;
assign i[3102]= 16'h1081;
assign i[3103]= 16'h103f;
assign i[3104]= 16'hfe1;
assign i[3105]= 16'hf74;
assign i[3106]= 16'hf04;
assign i[3107]= 16'hea1;
assign i[3108]= 16'he58;
assign i[3109]= 16'he36;
assign i[3110]= 16'he46;
assign i[3111]= 16'he92;
assign i[3112]= 16'hf21;
assign i[3113]= 16'hff8;
assign i[3114]= 16'h1119;
assign i[3115]= 16'h1284;
assign i[3116]= 16'h1434;
assign i[3117]= 16'h1622;
assign i[3118]= 16'h1846;
assign i[3119]= 16'h1a93;
assign i[3120]= 16'h1cfd;
assign i[3121]= 16'h1f73;
assign i[3122]= 16'h21e7;
assign i[3123]= 16'h2448;
assign i[3124]= 16'h2687;
assign i[3125]= 16'h2894;
assign i[3126]= 16'h2a65;
assign i[3127]= 16'h2bed;
assign i[3128]= 16'h2d25;
assign i[3129]= 16'h2e09;
assign i[3130]= 16'h2e98;
assign i[3131]= 16'h2ed4;
assign i[3132]= 16'h2ec4;
assign i[3133]= 16'h2e70;
assign i[3134]= 16'h2de5;
assign i[3135]= 16'h2d33;
assign i[3136]= 16'h2c69;
assign i[3137]= 16'h2b9b;
assign i[3138]= 16'h2ad9;
assign i[3139]= 16'h2a37;
assign i[3140]= 16'h29c4;
assign i[3141]= 16'h298f;
assign i[3142]= 16'h29a2;
assign i[3143]= 16'h2a05;
assign i[3144]= 16'h2aba;
assign i[3145]= 16'h2bbf;
assign i[3146]= 16'h2d0e;
assign i[3147]= 16'h2e99;
assign i[3148]= 16'h3050;
assign i[3149]= 16'h321e;
assign i[3150]= 16'h33e9;
assign i[3151]= 16'h3595;
assign i[3152]= 16'h3705;
assign i[3153]= 16'h381a;
assign i[3154]= 16'h38b7;
assign i[3155]= 16'h38be;
assign i[3156]= 16'h3818;
assign i[3157]= 16'h36b0;
assign i[3158]= 16'h3477;
assign i[3159]= 16'h3165;
assign i[3160]= 16'h2d79;
assign i[3161]= 16'h28bb;
assign i[3162]= 16'h2338;
assign i[3163]= 16'h1d08;
assign i[3164]= 16'h1649;
assign i[3165]= 16'hf20;
assign i[3166]= 16'h7b8;
assign i[3167]= 16'h40;
assign i[3168]= 16'hf8eb;
assign i[3169]= 16'hf1ea;
assign i[3170]= 16'heb72;
assign i[3171]= 16'he5b2;
assign i[3172]= 16'he0d6;
assign i[3173]= 16'hdd05;
assign i[3174]= 16'hda5e;
assign i[3175]= 16'hd8f7;
assign i[3176]= 16'hd8da;
assign i[3177]= 16'hda0b;
assign i[3178]= 16'hdc80;
assign i[3179]= 16'he024;
assign i[3180]= 16'he4da;
assign i[3181]= 16'hea79;
assign i[3182]= 16'hf0d1;
assign i[3183]= 16'hf7ad;
assign i[3184]= 16'hfed0;
assign i[3185]= 16'h5fc;
assign i[3186]= 16'hcf3;
assign i[3187]= 16'h1378;
assign i[3188]= 16'h1950;
assign i[3189]= 16'h1e49;
assign i[3190]= 16'h2236;
assign i[3191]= 16'h24f4;
assign i[3192]= 16'h266b;
assign i[3193]= 16'h268d;
assign i[3194]= 16'h255a;
assign i[3195]= 16'h22db;
assign i[3196]= 16'h1f28;
assign i[3197]= 16'h1a60;
assign i[3198]= 16'h14ac;
assign i[3199]= 16'he40;
assign i[3200]= 16'h752;
assign i[3201]= 16'h1d;
assign i[3202]= 16'hf8e1;
assign i[3203]= 16'hf1d6;
assign i[3204]= 16'heb39;
assign i[3205]= 16'he53f;
assign i[3206]= 16'he016;
assign i[3207]= 16'hdbe4;
assign i[3208]= 16'hd8c6;
assign i[3209]= 16'hd6d0;
assign i[3210]= 16'hd609;
assign i[3211]= 16'hd66e;
assign i[3212]= 16'hd7f2;
assign i[3213]= 16'hda7d;
assign i[3214]= 16'hddf1;
assign i[3215]= 16'he226;
assign i[3216]= 16'he6f0;
assign i[3217]= 16'hec1e;
assign i[3218]= 16'hf17e;
assign i[3219]= 16'hf6df;
assign i[3220]= 16'hfc0f;
assign i[3221]= 16'he2;
assign i[3222]= 16'h532;
assign i[3223]= 16'h8de;
assign i[3224]= 16'hbcc;
assign i[3225]= 16'hdec;
assign i[3226]= 16'hf35;
assign i[3227]= 16'hfa8;
assign i[3228]= 16'hf4d;
assign i[3229]= 16'he34;
assign i[3230]= 16'hc74;
assign i[3231]= 16'ha28;
assign i[3232]= 16'h771;
assign i[3233]= 16'h472;
assign i[3234]= 16'h14e;
assign i[3235]= 16'hfe2b;
assign i[3236]= 16'hfb2a;
assign i[3237]= 16'hf869;
assign i[3238]= 16'hf605;
assign i[3239]= 16'hf414;
assign i[3240]= 16'hf2a7;
assign i[3241]= 16'hf1c9;
assign i[3242]= 16'hf17f;
assign i[3243]= 16'hf1c7;
assign i[3244]= 16'hf29b;
assign i[3245]= 16'hf3f0;
assign i[3246]= 16'hf5b5;
assign i[3247]= 16'hf7d7;
assign i[3248]= 16'hfa3f;
assign i[3249]= 16'hfcd6;
assign i[3250]= 16'hff83;
assign i[3251]= 16'h22e;
assign i[3252]= 16'h4bf;
assign i[3253]= 16'h723;
assign i[3254]= 16'h945;
assign i[3255]= 16'hb16;
assign i[3256]= 16'hc89;
assign i[3257]= 16'hd95;
assign i[3258]= 16'he33;
assign i[3259]= 16'he61;
assign i[3260]= 16'he1f;
assign i[3261]= 16'hd6f;
assign i[3262]= 16'hc57;
assign i[3263]= 16'hadd;
assign i[3264]= 16'h90a;
assign i[3265]= 16'h6e7;
assign i[3266]= 16'h47d;
assign i[3267]= 16'h1d7;
assign i[3268]= 16'hff00;
assign i[3269]= 16'hfc00;
assign i[3270]= 16'hf8e1;
assign i[3271]= 16'hf5ae;
assign i[3272]= 16'hf26f;
assign i[3273]= 16'hef2d;
assign i[3274]= 16'hebf2;
assign i[3275]= 16'he8c6;
assign i[3276]= 16'he5b3;
assign i[3277]= 16'he2c1;
assign i[3278]= 16'hdffa;
assign i[3279]= 16'hdd67;
assign i[3280]= 16'hdb11;
assign i[3281]= 16'hd902;
assign i[3282]= 16'hd742;
assign i[3283]= 16'hd5d9;
assign i[3284]= 16'hd4cf;
assign i[3285]= 16'hd429;
assign i[3286]= 16'hd3ea;
assign i[3287]= 16'hd415;
assign i[3288]= 16'hd4a8;
assign i[3289]= 16'hd5a1;
assign i[3290]= 16'hd6f9;
assign i[3291]= 16'hd8a6;
assign i[3292]= 16'hda9d;
assign i[3293]= 16'hdcd0;
assign i[3294]= 16'hdf2c;
assign i[3295]= 16'he19f;
assign i[3296]= 16'he415;
assign i[3297]= 16'he679;
assign i[3298]= 16'he8b5;
assign i[3299]= 16'heab4;
assign i[3300]= 16'hec65;
assign i[3301]= 16'hedb6;
assign i[3302]= 16'hee9a;
assign i[3303]= 16'hef07;
assign i[3304]= 16'heef7;
assign i[3305]= 16'hee69;
assign i[3306]= 16'hed60;
assign i[3307]= 16'hebe5;
assign i[3308]= 16'hea04;
assign i[3309]= 16'he7d0;
assign i[3310]= 16'he55d;
assign i[3311]= 16'he2c3;
assign i[3312]= 16'he01e;
assign i[3313]= 16'hdd88;
assign i[3314]= 16'hdb1e;
assign i[3315]= 16'hd8fb;
assign i[3316]= 16'hd73a;
assign i[3317]= 16'hd5f1;
assign i[3318]= 16'hd533;
assign i[3319]= 16'hd510;
assign i[3320]= 16'hd591;
assign i[3321]= 16'hd6ba;
assign i[3322]= 16'hd88a;
assign i[3323]= 16'hdafa;
assign i[3324]= 16'hddfd;
assign i[3325]= 16'he181;
assign i[3326]= 16'he56f;
assign i[3327]= 16'he9ae;
assign i[3328]= 16'hee20;
assign i[3329]= 16'hf2a7;
assign i[3330]= 16'hf722;
assign i[3331]= 16'hfb73;
assign i[3332]= 16'hff7d;
assign i[3333]= 16'h323;
assign i[3334]= 16'h650;
assign i[3335]= 16'h8f0;
assign i[3336]= 16'haf4;
assign i[3337]= 16'hc54;
assign i[3338]= 16'hd0c;
assign i[3339]= 16'hd1f;
assign i[3340]= 16'hc94;
assign i[3341]= 16'hb79;
assign i[3342]= 16'h9df;
assign i[3343]= 16'h7da;
assign i[3344]= 16'h584;
assign i[3345]= 16'h2f5;
assign i[3346]= 16'h4a;
assign i[3347]= 16'hfd9d;
assign i[3348]= 16'hfb09;
assign i[3349]= 16'hf8a6;
assign i[3350]= 16'hf689;
assign i[3351]= 16'hf4c7;
assign i[3352]= 16'hf36e;
assign i[3353]= 16'hf288;
assign i[3354]= 16'hf21d;
assign i[3355]= 16'hf22f;
assign i[3356]= 16'hf2bb;
assign i[3357]= 16'hf3bd;
assign i[3358]= 16'hf52b;
assign i[3359]= 16'hf6f8;
assign i[3360]= 16'hf916;
assign i[3361]= 16'hfb74;
assign i[3362]= 16'hfe02;
assign i[3363]= 16'hac;
assign i[3364]= 16'h362;
assign i[3365]= 16'h612;
assign i[3366]= 16'h8ad;
assign i[3367]= 16'hb24;
assign i[3368]= 16'hd6c;
assign i[3369]= 16'hf79;
assign i[3370]= 16'h1145;
assign i[3371]= 16'h12ca;
assign i[3372]= 16'h1403;
assign i[3373]= 16'h14f0;
assign i[3374]= 16'h158f;
assign i[3375]= 16'h15e4;
assign i[3376]= 16'h15f0;
assign i[3377]= 16'h15b8;
assign i[3378]= 16'h153e;
assign i[3379]= 16'h1489;
assign i[3380]= 16'h139c;
assign i[3381]= 16'h127d;
assign i[3382]= 16'h1130;
assign i[3383]= 16'hfba;
assign i[3384]= 16'he21;
assign i[3385]= 16'hc68;
assign i[3386]= 16'ha94;
assign i[3387]= 16'h8aa;
assign i[3388]= 16'h6af;
assign i[3389]= 16'h4a9;
assign i[3390]= 16'h29d;
assign i[3391]= 16'h91;
assign i[3392]= 16'hfe8e;
assign i[3393]= 16'hfc97;
assign i[3394]= 16'hfab4;
assign i[3395]= 16'hf8ee;
assign i[3396]= 16'hf749;
assign i[3397]= 16'hf5ce;
assign i[3398]= 16'hf480;
assign i[3399]= 16'hf366;
assign i[3400]= 16'hf282;
assign i[3401]= 16'hf1d5;
assign i[3402]= 16'hf160;
assign i[3403]= 16'hf11f;
assign i[3404]= 16'hf110;
assign i[3405]= 16'hf12c;
assign i[3406]= 16'hf16a;
assign i[3407]= 16'hf1bf;
assign i[3408]= 16'hf222;
assign i[3409]= 16'hf284;
assign i[3410]= 16'hf2d9;
assign i[3411]= 16'hf313;
assign i[3412]= 16'hf324;
assign i[3413]= 16'hf302;
assign i[3414]= 16'hf2a1;
assign i[3415]= 16'hf1f8;
assign i[3416]= 16'hf103;
assign i[3417]= 16'hefbf;
assign i[3418]= 16'hee2c;
assign i[3419]= 16'hec4e;
assign i[3420]= 16'hea2e;
assign i[3421]= 16'he7d7;
assign i[3422]= 16'he556;
assign i[3423]= 16'he2bd;
assign i[3424]= 16'he01f;
assign i[3425]= 16'hdd90;
assign i[3426]= 16'hdb26;
assign i[3427]= 16'hd8f5;
assign i[3428]= 16'hd711;
assign i[3429]= 16'hd58c;
assign i[3430]= 16'hd476;
assign i[3431]= 16'hd3db;
assign i[3432]= 16'hd3c1;
assign i[3433]= 16'hd42b;
assign i[3434]= 16'hd519;
assign i[3435]= 16'hd683;
assign i[3436]= 16'hd85c;
assign i[3437]= 16'hda95;
assign i[3438]= 16'hdd1a;
assign i[3439]= 16'hdfd1;
assign i[3440]= 16'he2a2;
assign i[3441]= 16'he56f;
assign i[3442]= 16'he81c;
assign i[3443]= 16'hea8d;
assign i[3444]= 16'heca9;
assign i[3445]= 16'hee59;
assign i[3446]= 16'hef88;
assign i[3447]= 16'hf029;
assign i[3448]= 16'hf034;
assign i[3449]= 16'hefa5;
assign i[3450]= 16'hee81;
assign i[3451]= 16'hecd1;
assign i[3452]= 16'heaa5;
assign i[3453]= 16'he814;
assign i[3454]= 16'he538;
assign i[3455]= 16'he230;
assign i[3456]= 16'hdf1d;
assign i[3457]= 16'hdc22;
assign i[3458]= 16'hd963;
assign i[3459]= 16'hd700;
assign i[3460]= 16'hd51b;
assign i[3461]= 16'hd3ce;
assign i[3462]= 16'hd32f;
assign i[3463]= 16'hd34e;
assign i[3464]= 16'hd436;
assign i[3465]= 16'hd5e7;
assign i[3466]= 16'hd85c;
assign i[3467]= 16'hdb86;
assign i[3468]= 16'hdf53;
assign i[3469]= 16'he3a5;
assign i[3470]= 16'he85d;
assign i[3471]= 16'hed53;
assign i[3472]= 16'hf260;
assign i[3473]= 16'hf759;
assign i[3474]= 16'hfc13;
assign i[3475]= 16'h63;
assign i[3476]= 16'h426;
assign i[3477]= 16'h739;
assign i[3478]= 16'h981;
assign i[3479]= 16'hae7;
assign i[3480]= 16'hb60;
assign i[3481]= 16'hae6;
assign i[3482]= 16'h97f;
assign i[3483]= 16'h736;
assign i[3484]= 16'h41f;
assign i[3485]= 16'h59;
assign i[3486]= 16'hfc06;
assign i[3487]= 16'hf74c;
assign i[3488]= 16'hf258;
assign i[3489]= 16'hed58;
assign i[3490]= 16'he87b;
assign i[3491]= 16'he3ee;
assign i[3492]= 16'hdfda;
assign i[3493]= 16'hdc66;
assign i[3494]= 16'hd9b2;
assign i[3495]= 16'hd7d8;
assign i[3496]= 16'hd6e7;
assign i[3497]= 16'hd6e8;
assign i[3498]= 16'hd7dc;
assign i[3499]= 16'hd9b9;
assign i[3500]= 16'hdc6d;
assign i[3501]= 16'hdfdf;
assign i[3502]= 16'he3ef;
assign i[3503]= 16'he876;
assign i[3504]= 16'hed4b;
assign i[3505]= 16'hf240;
assign i[3506]= 16'hf729;
assign i[3507]= 16'hfbd7;
assign i[3508]= 16'h20;
assign i[3509]= 16'h3dd;
assign i[3510]= 16'h6ee;
assign i[3511]= 16'h934;
assign i[3512]= 16'ha9e;
assign i[3513]= 16'hb1f;
assign i[3514]= 16'hab2;
assign i[3515]= 16'h95d;
assign i[3516]= 16'h72b;
assign i[3517]= 16'h432;
assign i[3518]= 16'h8a;
assign i[3519]= 16'hfc57;
assign i[3520]= 16'hf7ba;
assign i[3521]= 16'hf2db;
assign i[3522]= 16'hede4;
assign i[3523]= 16'he8fe;
assign i[3524]= 16'he450;
assign i[3525]= 16'hdffe;
assign i[3526]= 16'hdc28;
assign i[3527]= 16'hd8eb;
assign i[3528]= 16'hd659;
assign i[3529]= 16'hd483;
assign i[3530]= 16'hd36e;
assign i[3531]= 16'hd31c;
assign i[3532]= 16'hd384;
assign i[3533]= 16'hd499;
assign i[3534]= 16'hd648;
assign i[3535]= 16'hd879;
assign i[3536]= 16'hdb0f;
assign i[3537]= 16'hddeb;
assign i[3538]= 16'he0ed;
assign i[3539]= 16'he3f4;
assign i[3540]= 16'he6df;
assign i[3541]= 16'he990;
assign i[3542]= 16'hebee;
assign i[3543]= 16'hede1;
assign i[3544]= 16'hef57;
assign i[3545]= 16'hf043;
assign i[3546]= 16'hf09e;
assign i[3547]= 16'hf067;
assign i[3548]= 16'hefa1;
assign i[3549]= 16'hee55;
assign i[3550]= 16'hec91;
assign i[3551]= 16'hea66;
assign i[3552]= 16'he7ea;
assign i[3553]= 16'he531;
assign i[3554]= 16'he254;
assign i[3555]= 16'hdf6c;
assign i[3556]= 16'hdc8f;
assign i[3557]= 16'hd9d3;
assign i[3558]= 16'hd74b;
assign i[3559]= 16'hd507;
assign i[3560]= 16'hd315;
assign i[3561]= 16'hd17b;
assign i[3562]= 16'hd040;
assign i[3563]= 16'hcf64;
assign i[3564]= 16'hcee3;
assign i[3565]= 16'hceb6;
assign i[3566]= 16'hced4;
assign i[3567]= 16'hcf31;
assign i[3568]= 16'hcfbe;
assign i[3569]= 16'hd06c;
assign i[3570]= 16'hd12b;
assign i[3571]= 16'hd1ec;
assign i[3572]= 16'hd2a2;
assign i[3573]= 16'hd341;
assign i[3574]= 16'hd3bd;
assign i[3575]= 16'hd411;
assign i[3576]= 16'hd436;
assign i[3577]= 16'hd42d;
assign i[3578]= 16'hd3f7;
assign i[3579]= 16'hd398;
assign i[3580]= 16'hd317;
assign i[3581]= 16'hd27e;
assign i[3582]= 16'hd1d9;
assign i[3583]= 16'hd133;
assign i[3584]= 16'hd09a;
assign i[3585]= 16'hd019;
assign i[3586]= 16'hcfbf;
assign i[3587]= 16'hcf95;
assign i[3588]= 16'hcfa5;
assign i[3589]= 16'hcff7;
assign i[3590]= 16'hd08f;
assign i[3591]= 16'hd16f;
assign i[3592]= 16'hd296;
assign i[3593]= 16'hd402;
assign i[3594]= 16'hd5ad;
assign i[3595]= 16'hd78d;
assign i[3596]= 16'hd99a;
assign i[3597]= 16'hdbc7;
assign i[3598]= 16'hde08;
assign i[3599]= 16'he04f;
assign i[3600]= 16'he290;
assign i[3601]= 16'he4bc;
assign i[3602]= 16'he6ca;
assign i[3603]= 16'he8ae;
assign i[3604]= 16'hea61;
assign i[3605]= 16'hebdc;
assign i[3606]= 16'hed1b;
assign i[3607]= 16'hee1d;
assign i[3608]= 16'heee2;
assign i[3609]= 16'hef6f;
assign i[3610]= 16'hefc8;
assign i[3611]= 16'heff4;
assign i[3612]= 16'heffd;
assign i[3613]= 16'hefec;
assign i[3614]= 16'hefcd;
assign i[3615]= 16'hefa9;
assign i[3616]= 16'hef8e;
assign i[3617]= 16'hef85;
assign i[3618]= 16'hef99;
assign i[3619]= 16'hefd4;
assign i[3620]= 16'hf03d;
assign i[3621]= 16'hf0db;
assign i[3622]= 16'hf1b5;
assign i[3623]= 16'hf2cf;
assign i[3624]= 16'hf42c;
assign i[3625]= 16'hf5cd;
assign i[3626]= 16'hf7b2;
assign i[3627]= 16'hf9dd;
assign i[3628]= 16'hfc49;
assign i[3629]= 16'hfef7;
assign i[3630]= 16'h1e0;
assign i[3631]= 16'h503;
assign i[3632]= 16'h85b;
assign i[3633]= 16'hbe2;
assign i[3634]= 16'hf91;
assign i[3635]= 16'h1363;
assign i[3636]= 16'h174f;
assign i[3637]= 16'h1b4d;
assign i[3638]= 16'h1f51;
assign i[3639]= 16'h2352;
assign i[3640]= 16'h2742;
assign i[3641]= 16'h2b14;
assign i[3642]= 16'h2eb8;
assign i[3643]= 16'h321f;
assign i[3644]= 16'h3537;
assign i[3645]= 16'h37ef;
assign i[3646]= 16'h3a34;
assign i[3647]= 16'h3bf6;
assign i[3648]= 16'h3d22;
assign i[3649]= 16'h3daa;
assign i[3650]= 16'h3d7f;
assign i[3651]= 16'h3c98;
assign i[3652]= 16'h3aeb;
assign i[3653]= 16'h3876;
assign i[3654]= 16'h3538;
assign i[3655]= 16'h3138;
assign i[3656]= 16'h2c7e;
assign i[3657]= 16'h271c;
assign i[3658]= 16'h2125;
assign i[3659]= 16'h1ab3;
assign i[3660]= 16'h13e4;
assign i[3661]= 16'hcdb;
assign i[3662]= 16'h5bc;
assign i[3663]= 16'hfeb0;
assign i[3664]= 16'hf7df;
assign i[3665]= 16'hf171;
assign i[3666]= 16'heb8e;
assign i[3667]= 16'he65c;
assign i[3668]= 16'he1fc;
assign i[3669]= 16'hde8a;
assign i[3670]= 16'hdc1e;
assign i[3671]= 16'hdac8;
assign i[3672]= 16'hda90;
assign i[3673]= 16'hdb78;
assign i[3674]= 16'hdd79;
assign i[3675]= 16'he083;
assign i[3676]= 16'he480;
assign i[3677]= 16'he952;
assign i[3678]= 16'heed5;
assign i[3679]= 16'hf4e1;
assign i[3680]= 16'hfb47;
assign i[3681]= 16'h1d9;
assign i[3682]= 16'h867;
assign i[3683]= 16'hec1;
assign i[3684]= 16'h14b8;
assign i[3685]= 16'h1a23;
assign i[3686]= 16'h1edb;
assign i[3687]= 16'h22c0;
assign i[3688]= 16'h25bb;
assign i[3689]= 16'h27ba;
assign i[3690]= 16'h28b3;
assign i[3691]= 16'h28a6;
assign i[3692]= 16'h2799;
assign i[3693]= 16'h259b;
assign i[3694]= 16'h22c2;
assign i[3695]= 16'h1f29;
assign i[3696]= 16'h1af0;
assign i[3697]= 16'h163c;
assign i[3698]= 16'h1133;
assign i[3699]= 16'hbfb;
assign i[3700]= 16'h6bd;
assign i[3701]= 16'h19c;
assign i[3702]= 16'hfcbd;
assign i[3703]= 16'hf83a;
assign i[3704]= 16'hf42e;
assign i[3705]= 16'hf0ac;
assign i[3706]= 16'hedc2;
assign i[3707]= 16'heb77;
assign i[3708]= 16'he9cc;
assign i[3709]= 16'he8bc;
assign i[3710]= 16'he83e;
assign i[3711]= 16'he843;
assign i[3712]= 16'he8b8;
assign i[3713]= 16'he98a;
assign i[3714]= 16'heaa1;
assign i[3715]= 16'hebe6;
assign i[3716]= 16'hed43;
assign i[3717]= 16'heea0;
assign i[3718]= 16'hefec;
assign i[3719]= 16'hf115;
assign i[3720]= 16'hf20e;
assign i[3721]= 16'hf2cf;
assign i[3722]= 16'hf351;
assign i[3723]= 16'hf393;
assign i[3724]= 16'hf398;
assign i[3725]= 16'hf366;
assign i[3726]= 16'hf306;
assign i[3727]= 16'hf284;
assign i[3728]= 16'hf1ee;
assign i[3729]= 16'hf152;
assign i[3730]= 16'hf0bf;
assign i[3731]= 16'hf044;
assign i[3732]= 16'hefee;
assign i[3733]= 16'hefca;
assign i[3734]= 16'hefe2;
assign i[3735]= 16'hf03d;
assign i[3736]= 16'hf0df;
assign i[3737]= 16'hf1cb;
assign i[3738]= 16'hf2ff;
assign i[3739]= 16'hf477;
assign i[3740]= 16'hf62c;
assign i[3741]= 16'hf815;
assign i[3742]= 16'hfa28;
assign i[3743]= 16'hfc57;
assign i[3744]= 16'hfe95;
assign i[3745]= 16'hd3;
assign i[3746]= 16'h305;
assign i[3747]= 16'h51b;
assign i[3748]= 16'h70a;
assign i[3749]= 16'h8c4;
assign i[3750]= 16'ha40;
assign i[3751]= 16'hb74;
assign i[3752]= 16'hc5a;
assign i[3753]= 16'hced;
assign i[3754]= 16'hd28;
assign i[3755]= 16'hd0a;
assign i[3756]= 16'hc93;
assign i[3757]= 16'hbc4;
assign i[3758]= 16'haa1;
assign i[3759]= 16'h92e;
assign i[3760]= 16'h76f;
assign i[3761]= 16'h56b;
assign i[3762]= 16'h327;
assign i[3763]= 16'had;
assign i[3764]= 16'hfe03;
assign i[3765]= 16'hfb30;
assign i[3766]= 16'hf83e;
assign i[3767]= 16'hf535;
assign i[3768]= 16'hf21e;
assign i[3769]= 16'hef02;
assign i[3770]= 16'hebeb;
assign i[3771]= 16'he8e2;
assign i[3772]= 16'he5f1;
assign i[3773]= 16'he321;
assign i[3774]= 16'he07d;
assign i[3775]= 16'hde0d;
assign i[3776]= 16'hdbdd;
assign i[3777]= 16'hd9f3;
assign i[3778]= 16'hd85a;
assign i[3779]= 16'hd718;
assign i[3780]= 16'hd636;
assign i[3781]= 16'hd5b8;
assign i[3782]= 16'hd5a3;
assign i[3783]= 16'hd5fa;
assign i[3784]= 16'hd6bf;
assign i[3785]= 16'hd7f3;
assign i[3786]= 16'hd992;
assign i[3787]= 16'hdb99;
assign i[3788]= 16'hde05;
assign i[3789]= 16'he0cc;
assign i[3790]= 16'he3e8;
assign i[3791]= 16'he74f;
assign i[3792]= 16'heaf6;
assign i[3793]= 16'heed1;
assign i[3794]= 16'hf2d4;
assign i[3795]= 16'hf6f3;
assign i[3796]= 16'hfb21;
assign i[3797]= 16'hff51;
assign i[3798]= 16'h377;
assign i[3799]= 16'h78a;
assign i[3800]= 16'hb7d;
assign i[3801]= 16'hf48;
assign i[3802]= 16'h12e2;
assign i[3803]= 16'h1646;
assign i[3804]= 16'h196c;
assign i[3805]= 16'h1c52;
assign i[3806]= 16'h1ef4;
assign i[3807]= 16'h2152;
assign i[3808]= 16'h236a;
assign i[3809]= 16'h253f;
assign i[3810]= 16'h26d3;
assign i[3811]= 16'h2827;
assign i[3812]= 16'h2941;
assign i[3813]= 16'h2a25;
assign i[3814]= 16'h2ad8;
assign i[3815]= 16'h2b5e;
assign i[3816]= 16'h2bbe;
assign i[3817]= 16'h2bfe;
assign i[3818]= 16'h2c23;
assign i[3819]= 16'h2c34;
assign i[3820]= 16'h2c35;
assign i[3821]= 16'h2c2c;
assign i[3822]= 16'h2c1f;
assign i[3823]= 16'h2c11;
assign i[3824]= 16'h2c08;
assign i[3825]= 16'h2c06;
assign i[3826]= 16'h2c0f;
assign i[3827]= 16'h2c25;
assign i[3828]= 16'h2c49;
assign i[3829]= 16'h2c7d;
assign i[3830]= 16'h2cbf;
assign i[3831]= 16'h2d10;
assign i[3832]= 16'h2d6d;
assign i[3833]= 16'h2dd3;
assign i[3834]= 16'h2e40;
assign i[3835]= 16'h2eaf;
assign i[3836]= 16'h2f1b;
assign i[3837]= 16'h2f80;
assign i[3838]= 16'h2fd7;
assign i[3839]= 16'h301b;
assign i[3840]= 16'h3046;
assign i[3841]= 16'h3053;
assign i[3842]= 16'h303c;
assign i[3843]= 16'h2ffe;
assign i[3844]= 16'h2f94;
assign i[3845]= 16'h2efc;
assign i[3846]= 16'h2e33;
assign i[3847]= 16'h2d3b;
assign i[3848]= 16'h2c12;
assign i[3849]= 16'h2abc;
assign i[3850]= 16'h293c;
assign i[3851]= 16'h2797;
assign i[3852]= 16'h25d2;
assign i[3853]= 16'h23f4;
assign i[3854]= 16'h2206;
assign i[3855]= 16'h200f;
assign i[3856]= 16'h1e1a;
assign i[3857]= 16'h1c2f;
assign i[3858]= 16'h1a57;
assign i[3859]= 16'h189d;
assign i[3860]= 16'h1708;
assign i[3861]= 16'h15a2;
assign i[3862]= 16'h1471;
assign i[3863]= 16'h137c;
assign i[3864]= 16'h12ca;
assign i[3865]= 16'h125e;
assign i[3866]= 16'h123b;
assign i[3867]= 16'h1264;
assign i[3868]= 16'h12da;
assign i[3869]= 16'h139b;
assign i[3870]= 16'h14a7;
assign i[3871]= 16'h15f9;
assign i[3872]= 16'h178f;
assign i[3873]= 16'h1962;
assign i[3874]= 16'h1b6c;
assign i[3875]= 16'h1da6;
assign i[3876]= 16'h2008;
assign i[3877]= 16'h2287;
assign i[3878]= 16'h251b;
assign i[3879]= 16'h27b7;
assign i[3880]= 16'h2a51;
assign i[3881]= 16'h2cdb;
assign i[3882]= 16'h2f49;
assign i[3883]= 16'h318d;
assign i[3884]= 16'h339b;
assign i[3885]= 16'h3563;
assign i[3886]= 16'h36da;
assign i[3887]= 16'h37f1;
assign i[3888]= 16'h389c;
assign i[3889]= 16'h38d2;
assign i[3890]= 16'h3886;
assign i[3891]= 16'h37b2;
assign i[3892]= 16'h364f;
assign i[3893]= 16'h3459;
assign i[3894]= 16'h31cf;
assign i[3895]= 16'h2eb2;
assign i[3896]= 16'h2b08;
assign i[3897]= 16'h26d8;
assign i[3898]= 16'h222c;
assign i[3899]= 16'h1d12;
assign i[3900]= 16'h179c;
assign i[3901]= 16'h11db;
assign i[3902]= 16'hbe7;
assign i[3903]= 16'h5d5;
assign i[3904]= 16'hffbf;
assign i[3905]= 16'hf9bd;
assign i[3906]= 16'hf3e8;
assign i[3907]= 16'hee59;
assign i[3908]= 16'he926;
assign i[3909]= 16'he466;
assign i[3910]= 16'he02b;
assign i[3911]= 16'hdc84;
assign i[3912]= 16'hd97d;
assign i[3913]= 16'hd720;
assign i[3914]= 16'hd570;
assign i[3915]= 16'hd46e;
assign i[3916]= 16'hd417;
assign i[3917]= 16'hd462;
assign i[3918]= 16'hd546;
assign i[3919]= 16'hd6b3;
assign i[3920]= 16'hd89a;
assign i[3921]= 16'hdae8;
assign i[3922]= 16'hdd8a;
assign i[3923]= 16'he06b;
assign i[3924]= 16'he377;
assign i[3925]= 16'he69a;
assign i[3926]= 16'he9c4;
assign i[3927]= 16'hece3;
assign i[3928]= 16'hefe9;
assign i[3929]= 16'hf2cc;
assign i[3930]= 16'hf584;
assign i[3931]= 16'hf80b;
assign i[3932]= 16'hfa5e;
assign i[3933]= 16'hfc7e;
assign i[3934]= 16'hfe6e;
assign i[3935]= 16'h32;
assign i[3936]= 16'h1d3;
assign i[3937]= 16'h357;
assign i[3938]= 16'h4c8;
assign i[3939]= 16'h62d;
assign i[3940]= 16'h791;
assign i[3941]= 16'h8fb;
assign i[3942]= 16'ha71;
assign i[3943]= 16'hbfa;
assign i[3944]= 16'hd99;
assign i[3945]= 16'hf50;
assign i[3946]= 16'h1121;
assign i[3947]= 16'h1309;
assign i[3948]= 16'h1506;
assign i[3949]= 16'h1713;
assign i[3950]= 16'h192c;
assign i[3951]= 16'h1b4a;
assign i[3952]= 16'h1d67;
assign i[3953]= 16'h1f7b;
assign i[3954]= 16'h2181;
assign i[3955]= 16'h2372;
assign i[3956]= 16'h254a;
assign i[3957]= 16'h2702;
assign i[3958]= 16'h2899;
assign i[3959]= 16'h2a0b;
assign i[3960]= 16'h2b56;
assign i[3961]= 16'h2c7b;
assign i[3962]= 16'h2d79;
assign i[3963]= 16'h2e50;
assign i[3964]= 16'h2f04;
assign i[3965]= 16'h2f94;
assign i[3966]= 16'h3004;
assign i[3967]= 16'h3054;
assign i[3968]= 16'h3087;
assign i[3969]= 16'h309d;
assign i[3970]= 16'h3099;
assign i[3971]= 16'h307b;
assign i[3972]= 16'h3044;
assign i[3973]= 16'h2ff4;
assign i[3974]= 16'h2f8e;
assign i[3975]= 16'h2f12;
assign i[3976]= 16'h2e82;
assign i[3977]= 16'h2de1;
assign i[3978]= 16'h2d32;
assign i[3979]= 16'h2c79;
assign i[3980]= 16'h2bbb;
assign i[3981]= 16'h2b00;
assign i[3982]= 16'h2a4d;
assign i[3983]= 16'h29ab;
assign i[3984]= 16'h2921;
assign i[3985]= 16'h28b9;
assign i[3986]= 16'h2879;
assign i[3987]= 16'h286a;
assign i[3988]= 16'h2892;
assign i[3989]= 16'h28f4;
assign i[3990]= 16'h2994;
assign i[3991]= 16'h2a71;
assign i[3992]= 16'h2b87;
assign i[3993]= 16'h2cd1;
assign i[3994]= 16'h2e45;
assign i[3995]= 16'h2fd6;
assign i[3996]= 16'h3176;
assign i[3997]= 16'h3311;
assign i[3998]= 16'h3493;
assign i[3999]= 16'h35e6;
assign i[4000]= 16'h36f3;
assign i[4001]= 16'h37a3;
assign i[4002]= 16'h37e0;
assign i[4003]= 16'h3794;
assign i[4004]= 16'h36af;
assign i[4005]= 16'h3522;
assign i[4006]= 16'h32e2;
assign i[4007]= 16'h2feb;
assign i[4008]= 16'h2c3d;
assign i[4009]= 16'h27df;
assign i[4010]= 16'h22dc;
assign i[4011]= 16'h1d48;
assign i[4012]= 16'h1738;
assign i[4013]= 16'h10ca;
assign i[4014]= 16'ha1f;
assign i[4015]= 16'h35a;
assign i[4016]= 16'hfca2;
assign i[4017]= 16'hf61d;
assign i[4018]= 16'heff1;
assign i[4019]= 16'hea44;
assign i[4020]= 16'he539;
assign i[4021]= 16'he0ec;
assign i[4022]= 16'hdd76;
assign i[4023]= 16'hdaea;
assign i[4024]= 16'hd954;
assign i[4025]= 16'hd8b8;
assign i[4026]= 16'hd914;
assign i[4027]= 16'hda5c;
assign i[4028]= 16'hdc80;
assign i[4029]= 16'hdf68;
assign i[4030]= 16'he2f6;
assign i[4031]= 16'he708;
assign i[4032]= 16'heb7a;
assign i[4033]= 16'hf022;
assign i[4034]= 16'hf4da;
assign i[4035]= 16'hf979;
assign i[4036]= 16'hfddb;
assign i[4037]= 16'h1db;
assign i[4038]= 16'h55e;
assign i[4039]= 16'h84b;
assign i[4040]= 16'ha8f;
assign i[4041]= 16'hc1f;
assign i[4042]= 16'hcf7;
assign i[4043]= 16'hd18;
assign i[4044]= 16'hc8c;
assign i[4045]= 16'hb62;
assign i[4046]= 16'h9af;
assign i[4047]= 16'h78d;
assign i[4048]= 16'h518;
assign i[4049]= 16'h270;
assign i[4050]= 16'hffb7;
assign i[4051]= 16'hfd0d;
assign i[4052]= 16'hfa91;
assign i[4053]= 16'hf863;
assign i[4054]= 16'hf69d;
assign i[4055]= 16'hf555;
assign i[4056]= 16'hf49e;
assign i[4057]= 16'hf486;
assign i[4058]= 16'hf514;
assign i[4059]= 16'hf64b;
assign i[4060]= 16'hf828;
assign i[4061]= 16'hfaa3;
assign i[4062]= 16'hfdb0;
assign i[4063]= 16'h13d;
assign i[4064]= 16'h53a;
assign i[4065]= 16'h98e;
assign i[4066]= 16'he21;
assign i[4067]= 16'h12dc;
assign i[4068]= 16'h17a4;
assign i[4069]= 16'h1c62;
assign i[4070]= 16'h20fd;
assign i[4071]= 16'h255f;
assign i[4072]= 16'h2975;
assign i[4073]= 16'h2d2e;
assign i[4074]= 16'h307c;
assign i[4075]= 16'h3352;
assign i[4076]= 16'h35a9;
assign i[4077]= 16'h377a;
assign i[4078]= 16'h38c2;
assign i[4079]= 16'h3980;
assign i[4080]= 16'h39b6;
assign i[4081]= 16'h3968;
assign i[4082]= 16'h389b;
assign i[4083]= 16'h3754;
assign i[4084]= 16'h359e;
assign i[4085]= 16'h337f;
assign i[4086]= 16'h3101;
assign i[4087]= 16'h2e2f;
assign i[4088]= 16'h2b14;
assign i[4089]= 16'h27b9;
assign i[4090]= 16'h242b;
assign i[4091]= 16'h2074;
assign i[4092]= 16'h1ca1;
assign i[4093]= 16'h18bd;
assign i[4094]= 16'h14d4;
assign i[4095]= 16'h10f2;
assign i[4096]= 16'hd23;
assign i[4097]= 16'h974;
assign i[4098]= 16'h5ef;
assign i[4099]= 16'h2a0;
assign i[4100]= 16'hff92;
assign i[4101]= 16'hfccf;
assign i[4102]= 16'hfa5f;
assign i[4103]= 16'hf84c;
assign i[4104]= 16'hf69c;
assign i[4105]= 16'hf554;
assign i[4106]= 16'hf478;
assign i[4107]= 16'hf40b;
assign i[4108]= 16'hf40d;
assign i[4109]= 16'hf47b;
assign i[4110]= 16'hf554;
assign i[4111]= 16'hf691;
assign i[4112]= 16'hf82c;
assign i[4113]= 16'hfa1c;
assign i[4114]= 16'hfc59;
assign i[4115]= 16'hfed7;
assign i[4116]= 16'h18a;
assign i[4117]= 16'h468;
assign i[4118]= 16'h765;
assign i[4119]= 16'ha73;
assign i[4120]= 16'hd87;
assign i[4121]= 16'h1097;
assign i[4122]= 16'h1396;
assign i[4123]= 16'h167d;
assign i[4124]= 16'h1943;
assign i[4125]= 16'h1be0;
assign i[4126]= 16'h1e4e;
assign i[4127]= 16'h2089;
assign i[4128]= 16'h228c;
assign i[4129]= 16'h2455;
assign i[4130]= 16'h25e2;
assign i[4131]= 16'h2732;
assign i[4132]= 16'h2845;
assign i[4133]= 16'h291c;
assign i[4134]= 16'h29b5;
assign i[4135]= 16'h2a14;
assign i[4136]= 16'h2a37;
assign i[4137]= 16'h2a21;
assign i[4138]= 16'h29d2;
assign i[4139]= 16'h294b;
assign i[4140]= 16'h288c;
assign i[4141]= 16'h2796;
assign i[4142]= 16'h2669;
assign i[4143]= 16'h2505;
assign i[4144]= 16'h236c;
assign i[4145]= 16'h219d;
assign i[4146]= 16'h1f98;
assign i[4147]= 16'h1d5f;
assign i[4148]= 16'h1af3;
assign i[4149]= 16'h1856;
assign i[4150]= 16'h1588;
assign i[4151]= 16'h128e;
assign i[4152]= 16'hf6a;
assign i[4153]= 16'hc1f;
assign i[4154]= 16'h8b1;
assign i[4155]= 16'h526;
assign i[4156]= 16'h181;
assign i[4157]= 16'hfdca;
assign i[4158]= 16'hfa05;
assign i[4159]= 16'hf637;
assign i[4160]= 16'hf268;
assign i[4161]= 16'hee9f;
assign i[4162]= 16'heae1;
assign i[4163]= 16'he735;
assign i[4164]= 16'he3a3;
assign i[4165]= 16'he031;
assign i[4166]= 16'hdce6;
assign i[4167]= 16'hd9c9;
assign i[4168]= 16'hd6e1;
assign i[4169]= 16'hd433;
assign i[4170]= 16'hd1c6;
assign i[4171]= 16'hcfa1;
assign i[4172]= 16'hcdc9;
assign i[4173]= 16'hcc44;
assign i[4174]= 16'hcb16;
assign i[4175]= 16'hca45;
assign i[4176]= 16'hc9d4;
assign i[4177]= 16'hc9c6;
assign i[4178]= 16'hca1d;
assign i[4179]= 16'hcada;
assign i[4180]= 16'hcbfd;
assign i[4181]= 16'hcd85;
assign i[4182]= 16'hcf6f;
assign i[4183]= 16'hd1b7;
assign i[4184]= 16'hd457;
assign i[4185]= 16'hd748;
assign i[4186]= 16'hda82;
assign i[4187]= 16'hddfa;
assign i[4188]= 16'he1a6;
assign i[4189]= 16'he578;
assign i[4190]= 16'he963;
assign i[4191]= 16'hed5a;
assign i[4192]= 16'hf14e;
assign i[4193]= 16'hf52e;
assign i[4194]= 16'hf8ee;
assign i[4195]= 16'hfc7d;
assign i[4196]= 16'hffcf;
assign i[4197]= 16'h2d4;
assign i[4198]= 16'h584;
assign i[4199]= 16'h7d4;
assign i[4200]= 16'h9b9;
assign i[4201]= 16'hb2f;
assign i[4202]= 16'hc30;
assign i[4203]= 16'hcb9;
assign i[4204]= 16'hccb;
assign i[4205]= 16'hc66;
assign i[4206]= 16'hb90;
assign i[4207]= 16'ha4c;
assign i[4208]= 16'h8a4;
assign i[4209]= 16'h6a0;
assign i[4210]= 16'h44b;
assign i[4211]= 16'h1af;
assign i[4212]= 16'hfedc;
assign i[4213]= 16'hfbdb;
assign i[4214]= 16'hf8ba;
assign i[4215]= 16'hf587;
assign i[4216]= 16'hf24f;
assign i[4217]= 16'hef1e;
assign i[4218]= 16'hebfe;
assign i[4219]= 16'he8fc;
assign i[4220]= 16'he61f;
assign i[4221]= 16'he371;
assign i[4222]= 16'he0f8;
assign i[4223]= 16'hdeb9;
assign i[4224]= 16'hdcba;
assign i[4225]= 16'hdafc;
assign i[4226]= 16'hd983;
assign i[4227]= 16'hd84d;
assign i[4228]= 16'hd75d;
assign i[4229]= 16'hd6af;
assign i[4230]= 16'hd643;
assign i[4231]= 16'hd616;
assign i[4232]= 16'hd625;
assign i[4233]= 16'hd66f;
assign i[4234]= 16'hd6ef;
assign i[4235]= 16'hd7a3;
assign i[4236]= 16'hd888;
assign i[4237]= 16'hd99c;
assign i[4238]= 16'hdadb;
assign i[4239]= 16'hdc43;
assign i[4240]= 16'hddd2;
assign i[4241]= 16'hdf86;
assign i[4242]= 16'he15d;
assign i[4243]= 16'he354;
assign i[4244]= 16'he56a;
assign i[4245]= 16'he79c;
assign i[4246]= 16'he9e6;
assign i[4247]= 16'hec47;
assign i[4248]= 16'heeba;
assign i[4249]= 16'hf13b;
assign i[4250]= 16'hf3c6;
assign i[4251]= 16'hf654;
assign i[4252]= 16'hf8e2;
assign i[4253]= 16'hfb67;
assign i[4254]= 16'hfddf;
assign i[4255]= 16'h41;
assign i[4256]= 16'h288;
assign i[4257]= 16'h4ad;
assign i[4258]= 16'h6a9;
assign i[4259]= 16'h878;
assign i[4260]= 16'ha13;
assign i[4261]= 16'hb78;
assign i[4262]= 16'hca4;
assign i[4263]= 16'hd95;
assign i[4264]= 16'he4c;
assign i[4265]= 16'heca;
assign i[4266]= 16'hf13;
assign i[4267]= 16'hf2d;
assign i[4268]= 16'hf1c;
assign i[4269]= 16'hee9;
assign i[4270]= 16'he9e;
assign i[4271]= 16'he42;
assign i[4272]= 16'hde1;
assign i[4273]= 16'hd84;
assign i[4274]= 16'hd34;
assign i[4275]= 16'hcfc;
assign i[4276]= 16'hce2;
assign i[4277]= 16'hced;
assign i[4278]= 16'hd21;
assign i[4279]= 16'hd80;
assign i[4280]= 16'he09;
assign i[4281]= 16'heba;
assign i[4282]= 16'hf8e;
assign i[4283]= 16'h107c;
assign i[4284]= 16'h117b;
assign i[4285]= 16'h127d;
assign i[4286]= 16'h1375;
assign i[4287]= 16'h1453;
assign i[4288]= 16'h1507;
assign i[4289]= 16'h1582;
assign i[4290]= 16'h15b4;
assign i[4291]= 16'h158e;
assign i[4292]= 16'h1505;
assign i[4293]= 16'h140d;
assign i[4294]= 16'h12a0;
assign i[4295]= 16'h10b9;
assign i[4296]= 16'he5a;
assign i[4297]= 16'hb85;
assign i[4298]= 16'h842;
assign i[4299]= 16'h49c;
assign i[4300]= 16'ha4;
assign i[4301]= 16'hfc6c;
assign i[4302]= 16'hf807;
assign i[4303]= 16'hf38f;
assign i[4304]= 16'hef1a;
assign i[4305]= 16'heac3;
assign i[4306]= 16'he6a3;
assign i[4307]= 16'he2d1;
assign i[4308]= 16'hdf62;
assign i[4309]= 16'hdc6b;
assign i[4310]= 16'hd9f9;
assign i[4311]= 16'hd81a;
assign i[4312]= 16'hd6d4;
assign i[4313]= 16'hd629;
assign i[4314]= 16'hd617;
assign i[4315]= 16'hd697;
assign i[4316]= 16'hd79c;
assign i[4317]= 16'hd918;
assign i[4318]= 16'hdaf5;
assign i[4319]= 16'hdd1e;
assign i[4320]= 16'hdf7a;
assign i[4321]= 16'he1ef;
assign i[4322]= 16'he464;
assign i[4323]= 16'he6bf;
assign i[4324]= 16'he8e7;
assign i[4325]= 16'heac8;
assign i[4326]= 16'hec50;
assign i[4327]= 16'hed6e;
assign i[4328]= 16'hee1a;
assign i[4329]= 16'hee4e;
assign i[4330]= 16'hee07;
assign i[4331]= 16'hed4a;
assign i[4332]= 16'hec1f;
assign i[4333]= 16'hea91;
assign i[4334]= 16'he8b2;
assign i[4335]= 16'he693;
assign i[4336]= 16'he44b;
assign i[4337]= 16'he1ef;
assign i[4338]= 16'hdf98;
assign i[4339]= 16'hdd5d;
assign i[4340]= 16'hdb56;
assign i[4341]= 16'hd998;
assign i[4342]= 16'hd836;
assign i[4343]= 16'hd741;
assign i[4344]= 16'hd6c7;
assign i[4345]= 16'hd6d2;
assign i[4346]= 16'hd768;
assign i[4347]= 16'hd88d;
assign i[4348]= 16'hda40;
assign i[4349]= 16'hdc7e;
assign i[4350]= 16'hdf40;
assign i[4351]= 16'he27b;
assign i[4352]= 16'he625;
assign i[4353]= 16'hea2f;
assign i[4354]= 16'hee8a;
assign i[4355]= 16'hf325;
assign i[4356]= 16'hf7f0;
assign i[4357]= 16'hfcd9;
assign i[4358]= 16'h1ce;
assign i[4359]= 16'h6c1;
assign i[4360]= 16'hba0;
assign i[4361]= 16'h105b;
assign i[4362]= 16'h14e4;
assign i[4363]= 16'h192d;
assign i[4364]= 16'h1d2a;
assign i[4365]= 16'h20cf;
assign i[4366]= 16'h2411;
assign i[4367]= 16'h26e8;
assign i[4368]= 16'h294a;
assign i[4369]= 16'h2b30;
assign i[4370]= 16'h2c96;
assign i[4371]= 16'h2d75;
assign i[4372]= 16'h2dcd;
assign i[4373]= 16'h2d9a;
assign i[4374]= 16'h2cde;
assign i[4375]= 16'h2b9c;
assign i[4376]= 16'h29d8;
assign i[4377]= 16'h2799;
assign i[4378]= 16'h24e9;
assign i[4379]= 16'h21d3;
assign i[4380]= 16'h1e66;
assign i[4381]= 16'h1ab1;
assign i[4382]= 16'h16c6;
assign i[4383]= 16'h12b9;
assign i[4384]= 16'he9f;
assign i[4385]= 16'ha8d;
assign i[4386]= 16'h699;
assign i[4387]= 16'h2d9;
assign i[4388]= 16'hff61;
assign i[4389]= 16'hfc43;
assign i[4390]= 16'hf990;
assign i[4391]= 16'hf756;
assign i[4392]= 16'hf5a0;
assign i[4393]= 16'hf476;
assign i[4394]= 16'hf3d9;
assign i[4395]= 16'hf3ca;
assign i[4396]= 16'hf444;
assign i[4397]= 16'hf53e;
assign i[4398]= 16'hf6ab;
assign i[4399]= 16'hf87e;
assign i[4400]= 16'hfaa3;
assign i[4401]= 16'hfd07;
assign i[4402]= 16'hff94;
assign i[4403]= 16'h235;
assign i[4404]= 16'h4d4;
assign i[4405]= 16'h75e;
assign i[4406]= 16'h9c0;
assign i[4407]= 16'hbea;
assign i[4408]= 16'hdce;
assign i[4409]= 16'hf64;
assign i[4410]= 16'h10a5;
assign i[4411]= 16'h118e;
assign i[4412]= 16'h1223;
assign i[4413]= 16'h1268;
assign i[4414]= 16'h1264;
assign i[4415]= 16'h1224;
assign i[4416]= 16'h11b4;
assign i[4417]= 16'h1123;
assign i[4418]= 16'h107f;
assign i[4419]= 16'hfd8;
assign i[4420]= 16'hf3b;
assign i[4421]= 16'heb6;
assign i[4422]= 16'he52;
assign i[4423]= 16'he17;
assign i[4424]= 16'he0b;
assign i[4425]= 16'he2d;
assign i[4426]= 16'he7d;
assign i[4427]= 16'hef4;
assign i[4428]= 16'hf8c;
assign i[4429]= 16'h1039;
assign i[4430]= 16'h10ee;
assign i[4431]= 16'h119d;
assign i[4432]= 16'h1237;
assign i[4433]= 16'h12aa;
assign i[4434]= 16'h12e9;
assign i[4435]= 16'h12e6;
assign i[4436]= 16'h1293;
assign i[4437]= 16'h11e7;
assign i[4438]= 16'h10da;
assign i[4439]= 16'hf69;
assign i[4440]= 16'hd90;
assign i[4441]= 16'hb53;
assign i[4442]= 16'h8b6;
assign i[4443]= 16'h5c1;
assign i[4444]= 16'h27e;
assign i[4445]= 16'hfefb;
assign i[4446]= 16'hfb44;
assign i[4447]= 16'hf76b;
assign i[4448]= 16'hf37e;
assign i[4449]= 16'hef8e;
assign i[4450]= 16'hebad;
assign i[4451]= 16'he7e9;
assign i[4452]= 16'he452;
assign i[4453]= 16'he0f4;
assign i[4454]= 16'hdddc;
assign i[4455]= 16'hdb16;
assign i[4456]= 16'hd8a9;
assign i[4457]= 16'hd69f;
assign i[4458]= 16'hd4fd;
assign i[4459]= 16'hd3c9;
assign i[4460]= 16'hd308;
assign i[4461]= 16'hd2bc;
assign i[4462]= 16'hd2e9;
assign i[4463]= 16'hd391;
assign i[4464]= 16'hd4b5;
assign i[4465]= 16'hd655;
assign i[4466]= 16'hd871;
assign i[4467]= 16'hdb08;
assign i[4468]= 16'hde17;
assign i[4469]= 16'he19b;
assign i[4470]= 16'he58d;
assign i[4471]= 16'he9e6;
assign i[4472]= 16'hee9a;
assign i[4473]= 16'hf39e;
assign i[4474]= 16'hf8e1;
assign i[4475]= 16'hfe52;
assign i[4476]= 16'h3da;
assign i[4477]= 16'h963;
assign i[4478]= 16'hed4;
assign i[4479]= 16'h1412;
assign i[4480]= 16'h1900;
assign i[4481]= 16'h1d83;
assign i[4482]= 16'h2180;
assign i[4483]= 16'h24de;
assign i[4484]= 16'h2786;
assign i[4485]= 16'h2966;
assign i[4486]= 16'h2a6f;
assign i[4487]= 16'h2a99;
assign i[4488]= 16'h29e2;
assign i[4489]= 16'h284d;
assign i[4490]= 16'h25e5;
assign i[4491]= 16'h22bc;
assign i[4492]= 16'h1eec;
assign i[4493]= 16'h1a91;
assign i[4494]= 16'h15d2;
assign i[4495]= 16'h10d5;
assign i[4496]= 16'hbc6;
assign i[4497]= 16'h6d2;
assign i[4498]= 16'h227;
assign i[4499]= 16'hfdef;
assign i[4500]= 16'hfa53;
assign i[4501]= 16'hf776;
assign i[4502]= 16'hf575;
assign i[4503]= 16'hf465;
assign i[4504]= 16'hf454;
assign i[4505]= 16'hf545;
assign i[4506]= 16'hf731;
assign i[4507]= 16'hfa0a;
assign i[4508]= 16'hfdb4;
assign i[4509]= 16'h20e;
assign i[4510]= 16'h6f0;
assign i[4511]= 16'hc29;
assign i[4512]= 16'h1184;
assign i[4513]= 16'h16cb;
assign i[4514]= 16'h1bc6;
assign i[4515]= 16'h2040;
assign i[4516]= 16'h2407;
assign i[4517]= 16'h26ed;
assign i[4518]= 16'h28cf;
assign i[4519]= 16'h298f;
assign i[4520]= 16'h291e;
assign i[4521]= 16'h2774;
assign i[4522]= 16'h2496;
assign i[4523]= 16'h2095;
assign i[4524]= 16'h1b8e;
assign i[4525]= 16'h15a6;
assign i[4526]= 16'hf0d;
assign i[4527]= 16'h7f9;
assign i[4528]= 16'ha6;
assign i[4529]= 16'hf954;
assign i[4530]= 16'hf240;
assign i[4531]= 16'hebab;
assign i[4532]= 16'he5cf;
assign i[4533]= 16'he0df;
assign i[4534]= 16'hdd09;
assign i[4535]= 16'hda6f;
assign i[4536]= 16'hd928;
assign i[4537]= 16'hd941;
assign i[4538]= 16'hdab8;
assign i[4539]= 16'hdd80;
assign i[4540]= 16'he17f;
assign i[4541]= 16'he692;
assign i[4542]= 16'hec8a;
assign i[4543]= 16'hf332;
assign i[4544]= 16'hfa4c;
assign i[4545]= 16'h199;
assign i[4546]= 16'h8d8;
assign i[4547]= 16'hfc7;
assign i[4548]= 16'h162a;
assign i[4549]= 16'h1bc6;
assign i[4550]= 16'h206d;
assign i[4551]= 16'h23f4;
assign i[4552]= 16'h263e;
assign i[4553]= 16'h2739;
assign i[4554]= 16'h26db;
assign i[4555]= 16'h252b;
assign i[4556]= 16'h2237;
assign i[4557]= 16'h1e19;
assign i[4558]= 16'h18f5;
assign i[4559]= 16'h12f5;
assign i[4560]= 16'hc4c;
assign i[4561]= 16'h52e;
assign i[4562]= 16'hfdd5;
assign i[4563]= 16'hf676;
assign i[4564]= 16'hef49;
assign i[4565]= 16'he881;
assign i[4566]= 16'he24b;
assign i[4567]= 16'hdcce;
assign i[4568]= 16'hd82a;
assign i[4569]= 16'hd475;
assign i[4570]= 16'hd1bd;
assign i[4571]= 16'hd007;
assign i[4572]= 16'hcf4f;
assign i[4573]= 16'hcf89;
assign i[4574]= 16'hd0a2;
assign i[4575]= 16'hd280;
assign i[4576]= 16'hd504;
assign i[4577]= 16'hd80d;
assign i[4578]= 16'hdb77;
assign i[4579]= 16'hdf1d;
assign i[4580]= 16'he2da;
assign i[4581]= 16'he68d;
assign i[4582]= 16'hea16;
assign i[4583]= 16'hed5c;
assign i[4584]= 16'hf047;
assign i[4585]= 16'hf2c9;
assign i[4586]= 16'hf4d4;
assign i[4587]= 16'hf664;
assign i[4588]= 16'hf779;
assign i[4589]= 16'hf816;
assign i[4590]= 16'hf845;
assign i[4591]= 16'hf812;
assign i[4592]= 16'hf78c;
assign i[4593]= 16'hf6c4;
assign i[4594]= 16'hf5cb;
assign i[4595]= 16'hf4b5;
assign i[4596]= 16'hf390;
assign i[4597]= 16'hf26f;
assign i[4598]= 16'hf15e;
assign i[4599]= 16'hf069;
assign i[4600]= 16'hef98;
assign i[4601]= 16'heef2;
assign i[4602]= 16'hee7a;
assign i[4603]= 16'hee30;
assign i[4604]= 16'hee12;
assign i[4605]= 16'hee1d;
assign i[4606]= 16'hee4a;
assign i[4607]= 16'hee93;
assign i[4608]= 16'heef0;
assign i[4609]= 16'hef5a;
assign i[4610]= 16'hefc9;
assign i[4611]= 16'hf036;
assign i[4612]= 16'hf09c;
assign i[4613]= 16'hf0f6;
assign i[4614]= 16'hf140;
assign i[4615]= 16'hf178;
assign i[4616]= 16'hf19e;
assign i[4617]= 16'hf1b2;
assign i[4618]= 16'hf1b6;
assign i[4619]= 16'hf1ad;
assign i[4620]= 16'hf198;
assign i[4621]= 16'hf17d;
assign i[4622]= 16'hf15e;
assign i[4623]= 16'hf13f;
assign i[4624]= 16'hf122;
assign i[4625]= 16'hf10a;
assign i[4626]= 16'hf0f8;
assign i[4627]= 16'hf0ed;
assign i[4628]= 16'hf0ea;
assign i[4629]= 16'hf0ec;
assign i[4630]= 16'hf0f4;
assign i[4631]= 16'hf0ff;
assign i[4632]= 16'hf10b;
assign i[4633]= 16'hf116;
assign i[4634]= 16'hf11d;
assign i[4635]= 16'hf120;
assign i[4636]= 16'hf11b;
assign i[4637]= 16'hf10f;
assign i[4638]= 16'hf0fc;
assign i[4639]= 16'hf0e1;
assign i[4640]= 16'hf0c0;
assign i[4641]= 16'hf09c;
assign i[4642]= 16'hf076;
assign i[4643]= 16'hf051;
assign i[4644]= 16'hf031;
assign i[4645]= 16'hf019;
assign i[4646]= 16'hf00a;
assign i[4647]= 16'hf009;
assign i[4648]= 16'hf016;
assign i[4649]= 16'hf032;
assign i[4650]= 16'hf05e;
assign i[4651]= 16'hf098;
assign i[4652]= 16'hf0df;
assign i[4653]= 16'hf12f;
assign i[4654]= 16'hf185;
assign i[4655]= 16'hf1db;
assign i[4656]= 16'hf22e;
assign i[4657]= 16'hf277;
assign i[4658]= 16'hf2b1;
assign i[4659]= 16'hf2d7;
assign i[4660]= 16'hf2e5;
assign i[4661]= 16'hf2d8;
assign i[4662]= 16'hf2ac;
assign i[4663]= 16'hf262;
assign i[4664]= 16'hf1fb;
assign i[4665]= 16'hf178;
assign i[4666]= 16'hf0de;
assign i[4667]= 16'hf032;
assign i[4668]= 16'hef7d;
assign i[4669]= 16'heec6;
assign i[4670]= 16'hee18;
assign i[4671]= 16'hed7c;
assign i[4672]= 16'hecfd;
assign i[4673]= 16'heca5;
assign i[4674]= 16'hec7e;
assign i[4675]= 16'hec90;
assign i[4676]= 16'hece3;
assign i[4677]= 16'hed7d;
assign i[4678]= 16'hee5f;
assign i[4679]= 16'hef8c;
assign i[4680]= 16'hf101;
assign i[4681]= 16'hf2bb;
assign i[4682]= 16'hf4b1;
assign i[4683]= 16'hf6db;
assign i[4684]= 16'hf92e;
assign i[4685]= 16'hfb9b;
assign i[4686]= 16'hfe14;
assign i[4687]= 16'h89;
assign i[4688]= 16'h2ea;
assign i[4689]= 16'h526;
assign i[4690]= 16'h72d;
assign i[4691]= 16'h8f2;
assign i[4692]= 16'ha66;
assign i[4693]= 16'hb7f;
assign i[4694]= 16'hc36;
assign i[4695]= 16'hc84;
assign i[4696]= 16'hc67;
assign i[4697]= 16'hbe2;
assign i[4698]= 16'haf7;
assign i[4699]= 16'h9b0;
assign i[4700]= 16'h818;
assign i[4701]= 16'h63b;
assign i[4702]= 16'h42a;
assign i[4703]= 16'h1f7;
assign i[4704]= 16'hffb8;
assign i[4705]= 16'hfd7e;
assign i[4706]= 16'hfb60;
assign i[4707]= 16'hf972;
assign i[4708]= 16'hf7c8;
assign i[4709]= 16'hf674;
assign i[4710]= 16'hf586;
assign i[4711]= 16'hf50c;
assign i[4712]= 16'hf510;
assign i[4713]= 16'hf599;
assign i[4714]= 16'hf6ad;
assign i[4715]= 16'hf84b;
assign i[4716]= 16'hfa6f;
assign i[4717]= 16'hfd14;
assign i[4718]= 16'h2d;
assign i[4719]= 16'h3af;
assign i[4720]= 16'h78a;
assign i[4721]= 16'hbac;
assign i[4722]= 16'h1000;
assign i[4723]= 16'h1472;
assign i[4724]= 16'h18eb;
assign i[4725]= 16'h1d57;
assign i[4726]= 16'h219f;
assign i[4727]= 16'h25b0;
assign i[4728]= 16'h2977;
assign i[4729]= 16'h2ce4;
assign i[4730]= 16'h2fe9;
assign i[4731]= 16'h327a;
assign i[4732]= 16'h3490;
assign i[4733]= 16'h3623;
assign i[4734]= 16'h3733;
assign i[4735]= 16'h37bf;
assign i[4736]= 16'h37cb;
assign i[4737]= 16'h375d;
assign i[4738]= 16'h367b;
assign i[4739]= 16'h3530;
assign i[4740]= 16'h3386;
assign i[4741]= 16'h3189;
assign i[4742]= 16'h2f44;
assign i[4743]= 16'h2cc3;
assign i[4744]= 16'h2a12;
assign i[4745]= 16'h273b;
assign i[4746]= 16'h2447;
assign i[4747]= 16'h213e;
assign i[4748]= 16'h1e26;
assign i[4749]= 16'h1b04;
assign i[4750]= 16'h17db;
assign i[4751]= 16'h14ae;
assign i[4752]= 16'h117d;
assign i[4753]= 16'he49;
assign i[4754]= 16'hb10;
assign i[4755]= 16'h7d4;
assign i[4756]= 16'h494;
assign i[4757]= 16'h151;
assign i[4758]= 16'hfe0e;
assign i[4759]= 16'hface;
assign i[4760]= 16'hf797;
assign i[4761]= 16'hf471;
assign i[4762]= 16'hf165;
assign i[4763]= 16'hee7f;
assign i[4764]= 16'hebcd;
assign i[4765]= 16'he95f;
assign i[4766]= 16'he743;
assign i[4767]= 16'he58b;
assign i[4768]= 16'he448;
assign i[4769]= 16'he389;
assign i[4770]= 16'he35c;
assign i[4771]= 16'he3cd;
assign i[4772]= 16'he4e5;
assign i[4773]= 16'he6a8;
assign i[4774]= 16'he919;
assign i[4775]= 16'hec31;
assign i[4776]= 16'hefe8;
assign i[4777]= 16'hf430;
assign i[4778]= 16'hf8f4;
assign i[4779]= 16'hfe1c;
assign i[4780]= 16'h389;
assign i[4781]= 16'h91d;
assign i[4782]= 16'heb2;
assign i[4783]= 16'h1421;
assign i[4784]= 16'h1945;
assign i[4785]= 16'h1df6;
assign i[4786]= 16'h2210;
assign i[4787]= 16'h2570;
assign i[4788]= 16'h27fa;
assign i[4789]= 16'h2994;
assign i[4790]= 16'h2a2d;
assign i[4791]= 16'h29b9;
assign i[4792]= 16'h2837;
assign i[4793]= 16'h25ab;
assign i[4794]= 16'h2223;
assign i[4795]= 16'h1db4;
assign i[4796]= 16'h187b;
assign i[4797]= 16'h129c;
assign i[4798]= 16'hc42;
assign i[4799]= 16'h599;
assign i[4800]= 16'hfed5;
assign i[4801]= 16'hf825;
assign i[4802]= 16'hf1bf;
assign i[4803]= 16'hebd2;
assign i[4804]= 16'he68d;
assign i[4805]= 16'he218;
assign i[4806]= 16'hde96;
assign i[4807]= 16'hdc22;
assign i[4808]= 16'hdad0;
assign i[4809]= 16'hdaaa;
assign i[4810]= 16'hdbb1;
assign i[4811]= 16'hdddd;
assign i[4812]= 16'he11d;
assign i[4813]= 16'he557;
assign i[4814]= 16'hea6d;
assign i[4815]= 16'hf037;
assign i[4816]= 16'hf68a;
assign i[4817]= 16'hfd37;
assign i[4818]= 16'h40e;
assign i[4819]= 16'hae0;
assign i[4820]= 16'h117e;
assign i[4821]= 16'h17ba;
assign i[4822]= 16'h1d70;
assign i[4823]= 16'h227b;
assign i[4824]= 16'h26c2;
assign i[4825]= 16'h2a30;
assign i[4826]= 16'h2cb8;
assign i[4827]= 16'h2e56;
assign i[4828]= 16'h2f0e;
assign i[4829]= 16'h2ee8;
assign i[4830]= 16'h2df5;
assign i[4831]= 16'h2c4c;
assign i[4832]= 16'h2a07;
assign i[4833]= 16'h2744;
assign i[4834]= 16'h2423;
assign i[4835]= 16'h20c6;
assign i[4836]= 16'h1d4e;
assign i[4837]= 16'h19d9;
assign i[4838]= 16'h1684;
assign i[4839]= 16'h1368;
assign i[4840]= 16'h109c;
assign i[4841]= 16'he2e;
assign i[4842]= 16'hc2a;
assign i[4843]= 16'ha97;
assign i[4844]= 16'h977;
assign i[4845]= 16'h8c5;
assign i[4846]= 16'h87a;
assign i[4847]= 16'h88c;
assign i[4848]= 16'h8eb;
assign i[4849]= 16'h988;
assign i[4850]= 16'ha51;
assign i[4851]= 16'hb33;
assign i[4852]= 16'hc1c;
assign i[4853]= 16'hcfa;
assign i[4854]= 16'hdbc;
assign i[4855]= 16'he56;
assign i[4856]= 16'heb9;
assign i[4857]= 16'hedc;
assign i[4858]= 16'heb8;
assign i[4859]= 16'he48;
assign i[4860]= 16'hd88;
assign i[4861]= 16'hc79;
assign i[4862]= 16'hb1d;
assign i[4863]= 16'h976;
assign i[4864]= 16'h78a;
assign i[4865]= 16'h55f;
assign i[4866]= 16'h2fa;
assign i[4867]= 16'h65;
assign i[4868]= 16'hfda6;
assign i[4869]= 16'hfac5;
assign i[4870]= 16'hf7c9;
assign i[4871]= 16'hf4bc;
assign i[4872]= 16'hf1a4;
assign i[4873]= 16'hee8a;
assign i[4874]= 16'heb76;
assign i[4875]= 16'he871;
assign i[4876]= 16'he583;
assign i[4877]= 16'he2b4;
assign i[4878]= 16'he00f;
assign i[4879]= 16'hdd9d;
assign i[4880]= 16'hdb67;
assign i[4881]= 16'hd977;
assign i[4882]= 16'hd7d7;
assign i[4883]= 16'hd690;
assign i[4884]= 16'hd5ac;
assign i[4885]= 16'hd531;
assign i[4886]= 16'hd527;
assign i[4887]= 16'hd593;
assign i[4888]= 16'hd677;
assign i[4889]= 16'hd7d5;
assign i[4890]= 16'hd9aa;
assign i[4891]= 16'hdbf3;
assign i[4892]= 16'hdea9;
assign i[4893]= 16'he1c2;
assign i[4894]= 16'he532;
assign i[4895]= 16'he8eb;
assign i[4896]= 16'hecdc;
assign i[4897]= 16'hf0f4;
assign i[4898]= 16'hf51f;
assign i[4899]= 16'hf94a;
assign i[4900]= 16'hfd61;
assign i[4901]= 16'h150;
assign i[4902]= 16'h508;
assign i[4903]= 16'h876;
assign i[4904]= 16'hb8e;
assign i[4905]= 16'he44;
assign i[4906]= 16'h1090;
assign i[4907]= 16'h126d;
assign i[4908]= 16'h13d9;
assign i[4909]= 16'h14d6;
assign i[4910]= 16'h1567;
assign i[4911]= 16'h1595;
assign i[4912]= 16'h1568;
assign i[4913]= 16'h14ed;
assign i[4914]= 16'h142e;
assign i[4915]= 16'h133b;
assign i[4916]= 16'h121f;
assign i[4917]= 16'h10e7;
assign i[4918]= 16'hfa0;
assign i[4919]= 16'he53;
assign i[4920]= 16'hd08;
assign i[4921]= 16'hbc5;
assign i[4922]= 16'ha8d;
assign i[4923]= 16'h960;
assign i[4924]= 16'h83c;
assign i[4925]= 16'h71c;
assign i[4926]= 16'h5fc;
assign i[4927]= 16'h4d1;
assign i[4928]= 16'h395;
assign i[4929]= 16'h23d;
assign i[4930]= 16'hbf;
assign i[4931]= 16'hff16;
assign i[4932]= 16'hfd36;
assign i[4933]= 16'hfb1d;
assign i[4934]= 16'hf8c7;
assign i[4935]= 16'hf635;
assign i[4936]= 16'hf369;
assign i[4937]= 16'hf06a;
assign i[4938]= 16'hed42;
assign i[4939]= 16'he9fc;
assign i[4940]= 16'he6a9;
assign i[4941]= 16'he35b;
assign i[4942]= 16'he025;
assign i[4943]= 16'hdd1e;
assign i[4944]= 16'hda5a;
assign i[4945]= 16'hd7f0;
assign i[4946]= 16'hd5f4;
assign i[4947]= 16'hd47c;
assign i[4948]= 16'hd397;
assign i[4949]= 16'hd354;
assign i[4950]= 16'hd3bf;
assign i[4951]= 16'hd4de;
assign i[4952]= 16'hd6b5;
assign i[4953]= 16'hd941;
assign i[4954]= 16'hdc7d;
assign i[4955]= 16'he05f;
assign i[4956]= 16'he4d9;
assign i[4957]= 16'he9d7;
assign i[4958]= 16'hef45;
assign i[4959]= 16'hf50b;
assign i[4960]= 16'hfb0e;
assign i[4961]= 16'h133;
assign i[4962]= 16'h75f;
assign i[4963]= 16'hd77;
assign i[4964]= 16'h135f;
assign i[4965]= 16'h18ff;
assign i[4966]= 16'h1e41;
assign i[4967]= 16'h2313;
assign i[4968]= 16'h2763;
assign i[4969]= 16'h2b26;
assign i[4970]= 16'h2e55;
assign i[4971]= 16'h30eb;
assign i[4972]= 16'h32ea;
assign i[4973]= 16'h3455;
assign i[4974]= 16'h3534;
assign i[4975]= 16'h3593;
assign i[4976]= 16'h357f;
assign i[4977]= 16'h3509;
assign i[4978]= 16'h3443;
assign i[4979]= 16'h333e;
assign i[4980]= 16'h320e;
assign i[4981]= 16'h30c6;
assign i[4982]= 16'h2f78;
assign i[4983]= 16'h2e33;
assign i[4984]= 16'h2d05;
assign i[4985]= 16'h2bfc;
assign i[4986]= 16'h2b1f;
assign i[4987]= 16'h2a76;
assign i[4988]= 16'h2a04;
assign i[4989]= 16'h29c9;
assign i[4990]= 16'h29c4;
assign i[4991]= 16'h29f1;
assign i[4992]= 16'h2a48;
assign i[4993]= 16'h2ac2;
assign i[4994]= 16'h2b56;
assign i[4995]= 16'h2bf8;
assign i[4996]= 16'h2c9f;
assign i[4997]= 16'h2d41;
assign i[4998]= 16'h2dd4;
assign i[4999]= 16'h2e51;
assign i[5000]= 16'h2eb0;
assign i[5001]= 16'h2eee;
assign i[5002]= 16'h2f07;
assign i[5003]= 16'h2efb;
assign i[5004]= 16'h2ecd;
assign i[5005]= 16'h2e7f;
assign i[5006]= 16'h2e17;
assign i[5007]= 16'h2d9d;
assign i[5008]= 16'h2d19;
assign i[5009]= 16'h2c94;
assign i[5010]= 16'h2c17;
assign i[5011]= 16'h2bab;
assign i[5012]= 16'h2b59;
assign i[5013]= 16'h2b27;
assign i[5014]= 16'h2b1b;
assign i[5015]= 16'h2b39;
assign i[5016]= 16'h2b82;
assign i[5017]= 16'h2bf4;
assign i[5018]= 16'h2c8c;
assign i[5019]= 16'h2d44;
assign i[5020]= 16'h2e13;
assign i[5021]= 16'h2eee;
assign i[5022]= 16'h2fca;
assign i[5023]= 16'h309a;
assign i[5024]= 16'h3150;
assign i[5025]= 16'h31df;
assign i[5026]= 16'h3238;
assign i[5027]= 16'h3251;
assign i[5028]= 16'h3220;
assign i[5029]= 16'h319c;
assign i[5030]= 16'h30c1;
assign i[5031]= 16'h2f8e;
assign i[5032]= 16'h2e03;
assign i[5033]= 16'h2c25;
assign i[5034]= 16'h29fe;
assign i[5035]= 16'h2799;
assign i[5036]= 16'h2504;
assign i[5037]= 16'h224f;
assign i[5038]= 16'h1f8f;
assign i[5039]= 16'h1cd6;
assign i[5040]= 16'h1a38;
assign i[5041]= 16'h17cb;
assign i[5042]= 16'h15a1;
assign i[5043]= 16'h13ca;
assign i[5044]= 16'h1257;
assign i[5045]= 16'h1152;
assign i[5046]= 16'h10c4;
assign i[5047]= 16'h10b1;
assign i[5048]= 16'h1118;
assign i[5049]= 16'h11f6;
assign i[5050]= 16'h1342;
assign i[5051]= 16'h14f0;
assign i[5052]= 16'h16ef;
assign i[5053]= 16'h192c;
assign i[5054]= 16'h1b93;
assign i[5055]= 16'h1e0c;
assign i[5056]= 16'h207f;
assign i[5057]= 16'h22d4;
assign i[5058]= 16'h24f3;
assign i[5059]= 16'h26c6;
assign i[5060]= 16'h283a;
assign i[5061]= 16'h293e;
assign i[5062]= 16'h29c5;
assign i[5063]= 16'h29c3;
assign i[5064]= 16'h2935;
assign i[5065]= 16'h2817;
assign i[5066]= 16'h266e;
assign i[5067]= 16'h243f;
assign i[5068]= 16'h2196;
assign i[5069]= 16'h1e80;
assign i[5070]= 16'h1b0e;
assign i[5071]= 16'h1754;
assign i[5072]= 16'h1366;
assign i[5073]= 16'hf5a;
assign i[5074]= 16'hb48;
assign i[5075]= 16'h745;
assign i[5076]= 16'h367;
assign i[5077]= 16'hffc3;
assign i[5078]= 16'hfc6a;
assign i[5079]= 16'hf96f;
assign i[5080]= 16'hf6dd;
assign i[5081]= 16'hf4c2;
assign i[5082]= 16'hf326;
assign i[5083]= 16'hf20f;
assign i[5084]= 16'hf180;
assign i[5085]= 16'hf179;
assign i[5086]= 16'hf1f9;
assign i[5087]= 16'hf2fc;
assign i[5088]= 16'hf47a;
assign i[5089]= 16'hf66b;
assign i[5090]= 16'hf8c6;
assign i[5091]= 16'hfb7f;
assign i[5092]= 16'hfe89;
assign i[5093]= 16'h1d6;
assign i[5094]= 16'h559;
assign i[5095]= 16'h903;
assign i[5096]= 16'hcc4;
assign i[5097]= 16'h108d;
assign i[5098]= 16'h144f;
assign i[5099]= 16'h17f9;
assign i[5100]= 16'h1b7e;
assign i[5101]= 16'h1ed0;
assign i[5102]= 16'h21e0;
assign i[5103]= 16'h24a2;
assign i[5104]= 16'h270c;
assign i[5105]= 16'h2914;
assign i[5106]= 16'h2ab1;
assign i[5107]= 16'h2bdf;
assign i[5108]= 16'h2c99;
assign i[5109]= 16'h2cdf;
assign i[5110]= 16'h2cb2;
assign i[5111]= 16'h2c16;
assign i[5112]= 16'h2b11;
assign i[5113]= 16'h29ae;
assign i[5114]= 16'h27f7;
assign i[5115]= 16'h25fa;
assign i[5116]= 16'h23c9;
assign i[5117]= 16'h2173;
assign i[5118]= 16'h1f0c;
assign i[5119]= 16'h1ca8;
assign i[5120]= 16'h1a59;
assign i[5121]= 16'h1832;
assign i[5122]= 16'h1646;
assign i[5123]= 16'h14a3;
assign i[5124]= 16'h1359;
assign i[5125]= 16'h1272;
assign i[5126]= 16'h11f5;
assign i[5127]= 16'h11e8;
assign i[5128]= 16'h124a;
assign i[5129]= 16'h1319;
assign i[5130]= 16'h144e;
assign i[5131]= 16'h15dc;
assign i[5132]= 16'h17b7;
assign i[5133]= 16'h19cd;
assign i[5134]= 16'h1c09;
assign i[5135]= 16'h1e57;
assign i[5136]= 16'h209e;
assign i[5137]= 16'h22c6;
assign i[5138]= 16'h24b9;
assign i[5139]= 16'h265e;
assign i[5140]= 16'h279f;
assign i[5141]= 16'h286b;
assign i[5142]= 16'h28af;
assign i[5143]= 16'h285d;
assign i[5144]= 16'h276d;
assign i[5145]= 16'h25d8;
assign i[5146]= 16'h239b;
assign i[5147]= 16'h20b8;
assign i[5148]= 16'h1d35;
assign i[5149]= 16'h191c;
assign i[5150]= 16'h147a;
assign i[5151]= 16'hf5e;
assign i[5152]= 16'h9dc;
assign i[5153]= 16'h409;
assign i[5154]= 16'hfdfc;
assign i[5155]= 16'hf7cc;
assign i[5156]= 16'hf191;
assign i[5157]= 16'heb64;
assign i[5158]= 16'he55d;
assign i[5159]= 16'hdf93;
assign i[5160]= 16'hda1d;
assign i[5161]= 16'hd50e;
assign i[5162]= 16'hd079;
assign i[5163]= 16'hcc6d;
assign i[5164]= 16'hc8fa;
assign i[5165]= 16'hc62a;
assign i[5166]= 16'hc405;
assign i[5167]= 16'hc293;
assign i[5168]= 16'hc1d5;
assign i[5169]= 16'hc1ce;
assign i[5170]= 16'hc279;
assign i[5171]= 16'hc3d4;
assign i[5172]= 16'hc5d5;
assign i[5173]= 16'hc873;
assign i[5174]= 16'hcba1;
assign i[5175]= 16'hcf50;
assign i[5176]= 16'hd36f;
assign i[5177]= 16'hd7e9;
assign i[5178]= 16'hdcaa;
assign i[5179]= 16'he19a;
assign i[5180]= 16'he6a2;
assign i[5181]= 16'heba9;
assign i[5182]= 16'hf095;
assign i[5183]= 16'hf54c;
assign i[5184]= 16'hf9b7;
assign i[5185]= 16'hfdbd;
assign i[5186]= 16'h148;
assign i[5187]= 16'h447;
assign i[5188]= 16'h6a8;
assign i[5189]= 16'h85d;
assign i[5190]= 16'h95e;
assign i[5191]= 16'h9a6;
assign i[5192]= 16'h933;
assign i[5193]= 16'h80c;
assign i[5194]= 16'h637;
assign i[5195]= 16'h3c4;
assign i[5196]= 16'hc4;
assign i[5197]= 16'hfd4f;
assign i[5198]= 16'hf97c;
assign i[5199]= 16'hf569;
assign i[5200]= 16'hf134;
assign i[5201]= 16'hecfe;
assign i[5202]= 16'he8e7;
assign i[5203]= 16'he50d;
assign i[5204]= 16'he191;
assign i[5205]= 16'hde8c;
assign i[5206]= 16'hdc16;
assign i[5207]= 16'hda45;
assign i[5208]= 16'hd927;
assign i[5209]= 16'hd8c6;
assign i[5210]= 16'hd926;
assign i[5211]= 16'hda45;
assign i[5212]= 16'hdc1d;
assign i[5213]= 16'hde9f;
assign i[5214]= 16'he1bb;
assign i[5215]= 16'he55a;
assign i[5216]= 16'he961;
assign i[5217]= 16'hedb3;
assign i[5218]= 16'hf231;
assign i[5219]= 16'hf6bb;
assign i[5220]= 16'hfb30;
assign i[5221]= 16'hff70;
assign i[5222]= 16'h35f;
assign i[5223]= 16'h6e3;
assign i[5224]= 16'h9e6;
assign i[5225]= 16'hc54;
assign i[5226]= 16'he20;
assign i[5227]= 16'hf42;
assign i[5228]= 16'hfb7;
assign i[5229]= 16'hf81;
assign i[5230]= 16'hea7;
assign i[5231]= 16'hd34;
assign i[5232]= 16'hb38;
assign i[5233]= 16'h8c5;
assign i[5234]= 16'h5f3;
assign i[5235]= 16'h2d7;
assign i[5236]= 16'hff8c;
assign i[5237]= 16'hfc29;
assign i[5238]= 16'hf8c7;
assign i[5239]= 16'hf57e;
assign i[5240]= 16'hf263;
assign i[5241]= 16'hef89;
assign i[5242]= 16'hed01;
assign i[5243]= 16'head7;
assign i[5244]= 16'he917;
assign i[5245]= 16'he7c7;
assign i[5246]= 16'he6eb;
assign i[5247]= 16'he684;
assign i[5248]= 16'he691;
assign i[5249]= 16'he70d;
assign i[5250]= 16'he7f2;
assign i[5251]= 16'he93a;
assign i[5252]= 16'headc;
assign i[5253]= 16'heccf;
assign i[5254]= 16'hef0a;
assign i[5255]= 16'hf183;
assign i[5256]= 16'hf433;
assign i[5257]= 16'hf710;
assign i[5258]= 16'hfa13;
assign i[5259]= 16'hfd35;
assign i[5260]= 16'h6f;
assign i[5261]= 16'h3bd;
assign i[5262]= 16'h71a;
assign i[5263]= 16'ha81;
assign i[5264]= 16'hded;
assign i[5265]= 16'h115a;
assign i[5266]= 16'h14c3;
assign i[5267]= 16'h1824;
assign i[5268]= 16'h1b76;
assign i[5269]= 16'h1eb4;
assign i[5270]= 16'h21d8;
assign i[5271]= 16'h24da;
assign i[5272]= 16'h27b2;
assign i[5273]= 16'h2a5a;
assign i[5274]= 16'h2cca;
assign i[5275]= 16'h2ef8;
assign i[5276]= 16'h30df;
assign i[5277]= 16'h3278;
assign i[5278]= 16'h33bc;
assign i[5279]= 16'h34a7;
assign i[5280]= 16'h3536;
assign i[5281]= 16'h3566;
assign i[5282]= 16'h3539;
assign i[5283]= 16'h34af;
assign i[5284]= 16'h33cd;
assign i[5285]= 16'h3298;
assign i[5286]= 16'h3118;
assign i[5287]= 16'h2f54;
assign i[5288]= 16'h2d58;
assign i[5289]= 16'h2b2f;
assign i[5290]= 16'h28e4;
assign i[5291]= 16'h2684;
assign i[5292]= 16'h241b;
assign i[5293]= 16'h21b6;
assign i[5294]= 16'h1f61;
assign i[5295]= 16'h1d25;
assign i[5296]= 16'h1b0d;
assign i[5297]= 16'h1920;
assign i[5298]= 16'h1764;
assign i[5299]= 16'h15df;
assign i[5300]= 16'h1492;
assign i[5301]= 16'h137f;
assign i[5302]= 16'h12a5;
assign i[5303]= 16'h1200;
assign i[5304]= 16'h118d;
assign i[5305]= 16'h1146;
assign i[5306]= 16'h1123;
assign i[5307]= 16'h111e;
assign i[5308]= 16'h112d;
assign i[5309]= 16'h1147;
assign i[5310]= 16'h1163;
assign i[5311]= 16'h1178;
assign i[5312]= 16'h117c;
assign i[5313]= 16'h1168;
assign i[5314]= 16'h1132;
assign i[5315]= 16'h10d4;
assign i[5316]= 16'h1046;
assign i[5317]= 16'hf82;
assign i[5318]= 16'he85;
assign i[5319]= 16'hd49;
assign i[5320]= 16'hbcc;
assign i[5321]= 16'ha0c;
assign i[5322]= 16'h808;
assign i[5323]= 16'h5c0;
assign i[5324]= 16'h336;
assign i[5325]= 16'h6a;
assign i[5326]= 16'hfd63;
assign i[5327]= 16'hfa22;
assign i[5328]= 16'hf6ae;
assign i[5329]= 16'hf30e;
assign i[5330]= 16'hef4a;
assign i[5331]= 16'heb6a;
assign i[5332]= 16'he779;
assign i[5333]= 16'he382;
assign i[5334]= 16'hdf91;
assign i[5335]= 16'hdbb4;
assign i[5336]= 16'hd7f8;
assign i[5337]= 16'hd46b;
assign i[5338]= 16'hd11d;
assign i[5339]= 16'hce1b;
assign i[5340]= 16'hcb73;
assign i[5341]= 16'hc935;
assign i[5342]= 16'hc76c;
assign i[5343]= 16'hc625;
assign i[5344]= 16'hc569;
assign i[5345]= 16'hc540;
assign i[5346]= 16'hc5b2;
assign i[5347]= 16'hc6c1;
assign i[5348]= 16'hc870;
assign i[5349]= 16'hcabb;
assign i[5350]= 16'hcda0;
assign i[5351]= 16'hd117;
assign i[5352]= 16'hd515;
assign i[5353]= 16'hd990;
assign i[5354]= 16'hde77;
assign i[5355]= 16'he3bb;
assign i[5356]= 16'he948;
assign i[5357]= 16'hef0a;
assign i[5358]= 16'hf4ec;
assign i[5359]= 16'hfada;
assign i[5360]= 16'hbb;
assign i[5361]= 16'h67d;
assign i[5362]= 16'hc0b;
assign i[5363]= 16'h1152;
assign i[5364]= 16'h163f;
assign i[5365]= 16'h1ac3;
assign i[5366]= 16'h1ed1;
assign i[5367]= 16'h225e;
assign i[5368]= 16'h2560;
assign i[5369]= 16'h27d2;
assign i[5370]= 16'h29b0;
assign i[5371]= 16'h2af8;
assign i[5372]= 16'h2bad;
assign i[5373]= 16'h2bd0;
assign i[5374]= 16'h2b68;
assign i[5375]= 16'h2a7c;
assign i[5376]= 16'h2913;
assign i[5377]= 16'h2739;
assign i[5378]= 16'h24f8;
assign i[5379]= 16'h225d;
assign i[5380]= 16'h1f73;
assign i[5381]= 16'h1c48;
assign i[5382]= 16'h18ea;
assign i[5383]= 16'h1567;
assign i[5384]= 16'h11cc;
assign i[5385]= 16'he27;
assign i[5386]= 16'ha87;
assign i[5387]= 16'h6f8;
assign i[5388]= 16'h389;
assign i[5389]= 16'h45;
assign i[5390]= 16'hfd3b;
assign i[5391]= 16'hfa75;
assign i[5392]= 16'hf7fd;
assign i[5393]= 16'hf5df;
assign i[5394]= 16'hf421;
assign i[5395]= 16'hf2cc;
assign i[5396]= 16'hf1e3;
assign i[5397]= 16'hf16c;
assign i[5398]= 16'hf165;
assign i[5399]= 16'hf1ce;
assign i[5400]= 16'hf2a3;
assign i[5401]= 16'hf3dd;
assign i[5402]= 16'hf572;
assign i[5403]= 16'hf758;
assign i[5404]= 16'hf97f;
assign i[5405]= 16'hfbd7;
assign i[5406]= 16'hfe4f;
assign i[5407]= 16'hd1;
assign i[5408]= 16'h34b;
assign i[5409]= 16'h5a8;
assign i[5410]= 16'h7d3;
assign i[5411]= 16'h9ba;
assign i[5412]= 16'hb4a;
assign i[5413]= 16'hc75;
assign i[5414]= 16'hd2f;
assign i[5415]= 16'hd70;
assign i[5416]= 16'hd33;
assign i[5417]= 16'hc79;
assign i[5418]= 16'hb46;
assign i[5419]= 16'h9a4;
assign i[5420]= 16'h7a1;
assign i[5421]= 16'h54f;
assign i[5422]= 16'h2c2;
assign i[5423]= 16'h15;
assign i[5424]= 16'hfd62;
assign i[5425]= 16'hfac4;
assign i[5426]= 16'hf859;
assign i[5427]= 16'hf63b;
assign i[5428]= 16'hf487;
assign i[5429]= 16'hf351;
assign i[5430]= 16'hf2af;
assign i[5431]= 16'hf2af;
assign i[5432]= 16'hf35b;
assign i[5433]= 16'hf4b7;
assign i[5434]= 16'hf6c1;
assign i[5435]= 16'hf970;
assign i[5436]= 16'hfcb7;
assign i[5437]= 16'h80;
assign i[5438]= 16'h4b5;
assign i[5439]= 16'h936;
assign i[5440]= 16'hde5;
assign i[5441]= 16'h129f;
assign i[5442]= 16'h1741;
assign i[5443]= 16'h1ba8;
assign i[5444]= 16'h1fb3;
assign i[5445]= 16'h2345;
assign i[5446]= 16'h2644;
assign i[5447]= 16'h289d;
assign i[5448]= 16'h2a40;
assign i[5449]= 16'h2b26;
assign i[5450]= 16'h2b50;
assign i[5451]= 16'h2ac3;
assign i[5452]= 16'h298d;
assign i[5453]= 16'h27c1;
assign i[5454]= 16'h2579;
assign i[5455]= 16'h22d3;
assign i[5456]= 16'h1ff0;
assign i[5457]= 16'h1cf4;
assign i[5458]= 16'h1a02;
assign i[5459]= 16'h173e;
assign i[5460]= 16'h14c9;
assign i[5461]= 16'h12c1;
assign i[5462]= 16'h113d;
assign i[5463]= 16'h1052;
assign i[5464]= 16'h100a;
assign i[5465]= 16'h106a;
assign i[5466]= 16'h116f;
assign i[5467]= 16'h130f;
assign i[5468]= 16'h1538;
assign i[5469]= 16'h17d2;
assign i[5470]= 16'h1abe;
assign i[5471]= 16'h1dd9;
assign i[5472]= 16'h20ff;
assign i[5473]= 16'h2407;
assign i[5474]= 16'h26c9;
assign i[5475]= 16'h291e;
assign i[5476]= 16'h2ae4;
assign i[5477]= 16'h2bfa;
assign i[5478]= 16'h2c47;
assign i[5479]= 16'h2bb8;
assign i[5480]= 16'h2a40;
assign i[5481]= 16'h27dd;
assign i[5482]= 16'h2493;
assign i[5483]= 16'h206e;
assign i[5484]= 16'h1b84;
assign i[5485]= 16'h15f0;
assign i[5486]= 16'hfd3;
assign i[5487]= 16'h956;
assign i[5488]= 16'h2a2;
assign i[5489]= 16'hfbe5;
assign i[5490]= 16'hf54c;
assign i[5491]= 16'hef03;
assign i[5492]= 16'he934;
assign i[5493]= 16'he407;
assign i[5494]= 16'hdf9c;
assign i[5495]= 16'hdc0e;
assign i[5496]= 16'hd972;
assign i[5497]= 16'hd7d5;
assign i[5498]= 16'hd73a;
assign i[5499]= 16'hd79f;
assign i[5500]= 16'hd8fb;
assign i[5501]= 16'hdb3a;
assign i[5502]= 16'hde45;
assign i[5503]= 16'he200;
assign i[5504]= 16'he649;
assign i[5505]= 16'heafc;
assign i[5506]= 16'heff4;
assign i[5507]= 16'hf50b;
assign i[5508]= 16'hfa1c;
assign i[5509]= 16'hff05;
assign i[5510]= 16'h3a6;
assign i[5511]= 16'h7e6;
assign i[5512]= 16'hbae;
assign i[5513]= 16'heee;
assign i[5514]= 16'h119b;
assign i[5515]= 16'h13b0;
assign i[5516]= 16'h152f;
assign i[5517]= 16'h161e;
assign i[5518]= 16'h1689;
assign i[5519]= 16'h167e;
assign i[5520]= 16'h1611;
assign i[5521]= 16'h1557;
assign i[5522]= 16'h1467;
assign i[5523]= 16'h135a;
assign i[5524]= 16'h1246;
assign i[5525]= 16'h1141;
assign i[5526]= 16'h1062;
assign i[5527]= 16'hfb8;
assign i[5528]= 16'hf54;
assign i[5529]= 16'hf40;
assign i[5530]= 16'hf86;
assign i[5531]= 16'h1028;
assign i[5532]= 16'h1127;
assign i[5533]= 16'h1281;
assign i[5534]= 16'h142f;
assign i[5535]= 16'h1627;
assign i[5536]= 16'h1860;
assign i[5537]= 16'h1aca;
assign i[5538]= 16'h1d59;
assign i[5539]= 16'h1ffd;
assign i[5540]= 16'h22a6;
assign i[5541]= 16'h2546;
assign i[5542]= 16'h27cf;
assign i[5543]= 16'h2a33;
assign i[5544]= 16'h2c68;
assign i[5545]= 16'h2e63;
assign i[5546]= 16'h301d;
assign i[5547]= 16'h318f;
assign i[5548]= 16'h32b5;
assign i[5549]= 16'h338d;
assign i[5550]= 16'h3415;
assign i[5551]= 16'h344f;
assign i[5552]= 16'h343a;
assign i[5553]= 16'h33da;
assign i[5554]= 16'h3332;
assign i[5555]= 16'h3246;
assign i[5556]= 16'h3118;
assign i[5557]= 16'h2fad;
assign i[5558]= 16'h2e07;
assign i[5559]= 16'h2c2b;
assign i[5560]= 16'h2a1a;
assign i[5561]= 16'h27d8;
assign i[5562]= 16'h2566;
assign i[5563]= 16'h22c6;
assign i[5564]= 16'h1ffb;
assign i[5565]= 16'h1d06;
assign i[5566]= 16'h19ea;
assign i[5567]= 16'h16a9;
assign i[5568]= 16'h1346;
assign i[5569]= 16'hfc7;
assign i[5570]= 16'hc2f;
assign i[5571]= 16'h885;
assign i[5572]= 16'h4d1;
assign i[5573]= 16'h11a;
assign i[5574]= 16'hfd6c;
assign i[5575]= 16'hf9cf;
assign i[5576]= 16'hf650;
assign i[5577]= 16'hf2fb;
assign i[5578]= 16'hefdf;
assign i[5579]= 16'hed08;
assign i[5580]= 16'hea83;
assign i[5581]= 16'he85e;
assign i[5582]= 16'he6a5;
assign i[5583]= 16'he562;
assign i[5584]= 16'he4a0;
assign i[5585]= 16'he467;
assign i[5586]= 16'he4ba;
assign i[5587]= 16'he59e;
assign i[5588]= 16'he713;
assign i[5589]= 16'he915;
assign i[5590]= 16'heb9f;
assign i[5591]= 16'heea8;
assign i[5592]= 16'hf223;
assign i[5593]= 16'hf603;
assign i[5594]= 16'hfa34;
assign i[5595]= 16'hfea4;
assign i[5596]= 16'h33b;
assign i[5597]= 16'h7e5;
assign i[5598]= 16'hc87;
assign i[5599]= 16'h1108;
assign i[5600]= 16'h1550;
assign i[5601]= 16'h1945;
assign i[5602]= 16'h1cd3;
assign i[5603]= 16'h1fe1;
assign i[5604]= 16'h225f;
assign i[5605]= 16'h243a;
assign i[5606]= 16'h2566;
assign i[5607]= 16'h25da;
assign i[5608]= 16'h258e;
assign i[5609]= 16'h2480;
assign i[5610]= 16'h22b3;
assign i[5611]= 16'h202a;
assign i[5612]= 16'h1cee;
assign i[5613]= 16'h190d;
assign i[5614]= 16'h1495;
assign i[5615]= 16'hf98;
assign i[5616]= 16'ha2b;
assign i[5617]= 16'h465;
assign i[5618]= 16'hfe5e;
assign i[5619]= 16'hf82d;
assign i[5620]= 16'hf1eb;
assign i[5621]= 16'hebb4;
assign i[5622]= 16'he59e;
assign i[5623]= 16'hdfc2;
assign i[5624]= 16'hda37;
assign i[5625]= 16'hd510;
assign i[5626]= 16'hd063;
assign i[5627]= 16'hcc3f;
assign i[5628]= 16'hc8b3;
assign i[5629]= 16'hc5cd;
assign i[5630]= 16'hc395;
assign i[5631]= 16'hc214;
assign i[5632]= 16'hc14e;
assign i[5633]= 16'hc146;
assign i[5634]= 16'hc1fc;
assign i[5635]= 16'hc36d;
assign i[5636]= 16'hc593;
assign i[5637]= 16'hc869;
assign i[5638]= 16'hcbe2;
assign i[5639]= 16'hcff5;
assign i[5640]= 16'hd492;
assign i[5641]= 16'hd9a8;
assign i[5642]= 16'hdf27;
assign i[5643]= 16'he4fa;
assign i[5644]= 16'heb0b;
assign i[5645]= 16'hf145;
assign i[5646]= 16'hf78f;
assign i[5647]= 16'hfdd1;
assign i[5648]= 16'h3f3;
assign i[5649]= 16'h9de;
assign i[5650]= 16'hf7c;
assign i[5651]= 16'h14b5;
assign i[5652]= 16'h1976;
assign i[5653]= 16'h1dae;
assign i[5654]= 16'h214e;
assign i[5655]= 16'h244a;
assign i[5656]= 16'h269c;
assign i[5657]= 16'h2840;
assign i[5658]= 16'h2935;
assign i[5659]= 16'h2982;
assign i[5660]= 16'h292e;
assign i[5661]= 16'h2848;
assign i[5662]= 16'h26de;
assign i[5663]= 16'h2507;
assign i[5664]= 16'h22d7;
assign i[5665]= 16'h2068;
assign i[5666]= 16'h1dd3;
assign i[5667]= 16'h1b32;
assign i[5668]= 16'h189d;
assign i[5669]= 16'h162d;
assign i[5670]= 16'h13f5;
assign i[5671]= 16'h1209;
assign i[5672]= 16'h1076;
assign i[5673]= 16'hf45;
assign i[5674]= 16'he79;
assign i[5675]= 16'he13;
assign i[5676]= 16'he0c;
assign i[5677]= 16'he59;
assign i[5678]= 16'heea;
assign i[5679]= 16'hfaa;
assign i[5680]= 16'h1084;
assign i[5681]= 16'h115e;
assign i[5682]= 16'h121c;
assign i[5683]= 16'h12a5;
assign i[5684]= 16'h12df;
assign i[5685]= 16'h12b3;
assign i[5686]= 16'h120c;
assign i[5687]= 16'h10dc;
assign i[5688]= 16'hf18;
assign i[5689]= 16'hcbb;
assign i[5690]= 16'h9c8;
assign i[5691]= 16'h648;
assign i[5692]= 16'h249;
assign i[5693]= 16'hfde1;
assign i[5694]= 16'hf928;
assign i[5695]= 16'hf43f;
assign i[5696]= 16'hef48;
assign i[5697]= 16'hea67;
assign i[5698]= 16'he5c3;
assign i[5699]= 16'he180;
assign i[5700]= 16'hddc1;
assign i[5701]= 16'hdaa5;
assign i[5702]= 16'hd849;
assign i[5703]= 16'hd6c0;
assign i[5704]= 16'hd619;
assign i[5705]= 16'hd65a;
assign i[5706]= 16'hd783;
assign i[5707]= 16'hd98a;
assign i[5708]= 16'hdc5e;
assign i[5709]= 16'hdfe9;
assign i[5710]= 16'he40a;
assign i[5711]= 16'he8a0;
assign i[5712]= 16'hed82;
assign i[5713]= 16'hf287;
assign i[5714]= 16'hf784;
assign i[5715]= 16'hfc4e;
assign i[5716]= 16'hbd;
assign i[5717]= 16'h4af;
assign i[5718]= 16'h804;
assign i[5719]= 16'haa5;
assign i[5720]= 16'hc7f;
assign i[5721]= 16'hd8b;
assign i[5722]= 16'hdc7;
assign i[5723]= 16'hd3b;
assign i[5724]= 16'hbf7;
assign i[5725]= 16'ha10;
assign i[5726]= 16'h7a5;
assign i[5727]= 16'h4d6;
assign i[5728]= 16'h1cb;
assign i[5729]= 16'hfeac;
assign i[5730]= 16'hfba0;
assign i[5731]= 16'hf8d0;
assign i[5732]= 16'hf661;
assign i[5733]= 16'hf474;
assign i[5734]= 16'hf324;
assign i[5735]= 16'hf288;
assign i[5736]= 16'hf2ae;
assign i[5737]= 16'hf39c;
assign i[5738]= 16'hf552;
assign i[5739]= 16'hf7c7;
assign i[5740]= 16'hfaea;
assign i[5741]= 16'hfea6;
assign i[5742]= 16'h2dc;
assign i[5743]= 16'h76e;
assign i[5744]= 16'hc37;
assign i[5745]= 16'h1113;
assign i[5746]= 16'h15db;
assign i[5747]= 16'h1a6a;
assign i[5748]= 16'h1ea0;
assign i[5749]= 16'h225d;
assign i[5750]= 16'h2589;
assign i[5751]= 16'h2811;
assign i[5752]= 16'h29e7;
assign i[5753]= 16'h2b05;
assign i[5754]= 16'h2b6c;
assign i[5755]= 16'h2b23;
assign i[5756]= 16'h2a37;
assign i[5757]= 16'h28bb;
assign i[5758]= 16'h26c6;
assign i[5759]= 16'h2473;
assign i[5760]= 16'h21e0;
assign i[5761]= 16'h1f2b;
assign i[5762]= 16'h1c73;
assign i[5763]= 16'h19d6;
assign i[5764]= 16'h176f;
assign i[5765]= 16'h1557;
assign i[5766]= 16'h13a2;
assign i[5767]= 16'h125f;
assign i[5768]= 16'h119b;
assign i[5769]= 16'h1159;
assign i[5770]= 16'h119a;
assign i[5771]= 16'h125a;
assign i[5772]= 16'h138e;
assign i[5773]= 16'h1528;
assign i[5774]= 16'h1716;
assign i[5775]= 16'h1944;
assign i[5776]= 16'h1b9b;
assign i[5777]= 16'h1e02;
assign i[5778]= 16'h2061;
assign i[5779]= 16'h229f;
assign i[5780]= 16'h24a6;
assign i[5781]= 16'h2660;
assign i[5782]= 16'h27bb;
assign i[5783]= 16'h28a5;
assign i[5784]= 16'h2914;
assign i[5785]= 16'h28fc;
assign i[5786]= 16'h2858;
assign i[5787]= 16'h2727;
assign i[5788]= 16'h2569;
assign i[5789]= 16'h2322;
assign i[5790]= 16'h205b;
assign i[5791]= 16'h1d1c;
assign i[5792]= 16'h1973;
assign i[5793]= 16'h156d;
assign i[5794]= 16'h111a;
assign i[5795]= 16'hc8b;
assign i[5796]= 16'h7d0;
assign i[5797]= 16'h2fb;
assign i[5798]= 16'hfe1e;
assign i[5799]= 16'hf949;
assign i[5800]= 16'hf48c;
assign i[5801]= 16'heff7;
assign i[5802]= 16'heb98;
assign i[5803]= 16'he77c;
assign i[5804]= 16'he3af;
assign i[5805]= 16'he03b;
assign i[5806]= 16'hdd28;
assign i[5807]= 16'hda7d;
assign i[5808]= 16'hd83e;
assign i[5809]= 16'hd670;
assign i[5810]= 16'hd513;
assign i[5811]= 16'hd426;
assign i[5812]= 16'hd3a8;
assign i[5813]= 16'hd394;
assign i[5814]= 16'hd3e4;
assign i[5815]= 16'hd491;
assign i[5816]= 16'hd592;
assign i[5817]= 16'hd6dd;
assign i[5818]= 16'hd867;
assign i[5819]= 16'hda23;
assign i[5820]= 16'hdc04;
assign i[5821]= 16'hddfe;
assign i[5822]= 16'he002;
assign i[5823]= 16'he203;
assign i[5824]= 16'he3f6;
assign i[5825]= 16'he5cd;
assign i[5826]= 16'he77d;
assign i[5827]= 16'he8fd;
assign i[5828]= 16'hea44;
assign i[5829]= 16'heb4b;
assign i[5830]= 16'hec0c;
assign i[5831]= 16'hec85;
assign i[5832]= 16'hecb4;
assign i[5833]= 16'hec98;
assign i[5834]= 16'hec33;
assign i[5835]= 16'heb89;
assign i[5836]= 16'hea9e;
assign i[5837]= 16'he979;
assign i[5838]= 16'he820;
assign i[5839]= 16'he69c;
assign i[5840]= 16'he4f6;
assign i[5841]= 16'he336;
assign i[5842]= 16'he169;
assign i[5843]= 16'hdf96;
assign i[5844]= 16'hddc9;
assign i[5845]= 16'hdc0c;
assign i[5846]= 16'hda69;
assign i[5847]= 16'hd8ea;
assign i[5848]= 16'hd798;
assign i[5849]= 16'hd67d;
assign i[5850]= 16'hd5a1;
assign i[5851]= 16'hd50d;
assign i[5852]= 16'hd4c7;
assign i[5853]= 16'hd4d7;
assign i[5854]= 16'hd542;
assign i[5855]= 16'hd60c;
assign i[5856]= 16'hd739;
assign i[5857]= 16'hd8cb;
assign i[5858]= 16'hdac2;
assign i[5859]= 16'hdd1b;
assign i[5860]= 16'hdfd3;
assign i[5861]= 16'he2e5;
assign i[5862]= 16'he646;
assign i[5863]= 16'he9ed;
assign i[5864]= 16'hedcd;
assign i[5865]= 16'hf1d6;
assign i[5866]= 16'hf5f5;
assign i[5867]= 16'hfa18;
assign i[5868]= 16'hfe2a;
assign i[5869]= 16'h212;
assign i[5870]= 16'h5bc;
assign i[5871]= 16'h910;
assign i[5872]= 16'hbf8;
assign i[5873]= 16'he5f;
assign i[5874]= 16'h1032;
assign i[5875]= 16'h1162;
assign i[5876]= 16'h11e1;
assign i[5877]= 16'h11a9;
assign i[5878]= 16'h10b4;
assign i[5879]= 16'hf05;
assign i[5880]= 16'hca3;
assign i[5881]= 16'h999;
assign i[5882]= 16'h5fa;
assign i[5883]= 16'h1db;
assign i[5884]= 16'hfd5a;
assign i[5885]= 16'hf892;
assign i[5886]= 16'hf3a8;
assign i[5887]= 16'heec0;
assign i[5888]= 16'hea01;
assign i[5889]= 16'he58f;
assign i[5890]= 16'he190;
assign i[5891]= 16'hde25;
assign i[5892]= 16'hdb6f;
assign i[5893]= 16'hd986;
assign i[5894]= 16'hd880;
assign i[5895]= 16'hd86c;
assign i[5896]= 16'hd94f;
assign i[5897]= 16'hdb2c;
assign i[5898]= 16'hddf9;
assign i[5899]= 16'he1a9;
assign i[5900]= 16'he624;
assign i[5901]= 16'heb4f;
assign i[5902]= 16'hf107;
assign i[5903]= 16'hf725;
assign i[5904]= 16'hfd7e;
assign i[5905]= 16'h3e5;
assign i[5906]= 16'ha2c;
assign i[5907]= 16'h1025;
assign i[5908]= 16'h15a5;
assign i[5909]= 16'h1a82;
assign i[5910]= 16'h1e99;
assign i[5911]= 16'h21cb;
assign i[5912]= 16'h23fe;
assign i[5913]= 16'h2521;
assign i[5914]= 16'h252b;
assign i[5915]= 16'h2419;
assign i[5916]= 16'h21ef;
assign i[5917]= 16'h1ebb;
assign i[5918]= 16'h1a91;
assign i[5919]= 16'h1589;
assign i[5920]= 16'hfc3;
assign i[5921]= 16'h963;
assign i[5922]= 16'h28e;
assign i[5923]= 16'hfb6e;
assign i[5924]= 16'hf42a;
assign i[5925]= 16'hecec;
assign i[5926]= 16'he5db;
assign i[5927]= 16'hdf1c;
assign i[5928]= 16'hd8d1;
assign i[5929]= 16'hd317;
assign i[5930]= 16'hce07;
assign i[5931]= 16'hc9b4;
assign i[5932]= 16'hc62c;
assign i[5933]= 16'hc37a;
assign i[5934]= 16'hc1a0;
assign i[5935]= 16'hc09f;
assign i[5936]= 16'hc071;
assign i[5937]= 16'hc10e;
assign i[5938]= 16'hc269;
assign i[5939]= 16'hc475;
assign i[5940]= 16'hc720;
assign i[5941]= 16'hca59;
assign i[5942]= 16'hce0d;
assign i[5943]= 16'hd22c;
assign i[5944]= 16'hd6a2;
assign i[5945]= 16'hdb5f;
assign i[5946]= 16'he053;
assign i[5947]= 16'he570;
assign i[5948]= 16'heaa9;
assign i[5949]= 16'heff3;
assign i[5950]= 16'hf542;
assign i[5951]= 16'hfa90;
assign i[5952]= 16'hffd2;
assign i[5953]= 16'h502;
assign i[5954]= 16'ha1b;
assign i[5955]= 16'hf16;
assign i[5956]= 16'h13ec;
assign i[5957]= 16'h1896;
assign i[5958]= 16'h1d0f;
assign i[5959]= 16'h214f;
assign i[5960]= 16'h254f;
assign i[5961]= 16'h2905;
assign i[5962]= 16'h2c6b;
assign i[5963]= 16'h2f78;
assign i[5964]= 16'h3222;
assign i[5965]= 16'h3462;
assign i[5966]= 16'h3631;
assign i[5967]= 16'h3787;
assign i[5968]= 16'h385e;
assign i[5969]= 16'h38b3;
assign i[5970]= 16'h3883;
assign i[5971]= 16'h37cd;
assign i[5972]= 16'h3693;
assign i[5973]= 16'h34d8;
assign i[5974]= 16'h32a3;
assign i[5975]= 16'h2ffb;
assign i[5976]= 16'h2ceb;
assign i[5977]= 16'h297e;
assign i[5978]= 16'h25c4;
assign i[5979]= 16'h21cb;
assign i[5980]= 16'h1da5;
assign i[5981]= 16'h1962;
assign i[5982]= 16'h1516;
assign i[5983]= 16'h10d1;
assign i[5984]= 16'hca6;
assign i[5985]= 16'h8a6;
assign i[5986]= 16'h4e0;
assign i[5987]= 16'h164;
assign i[5988]= 16'hfe3f;
assign i[5989]= 16'hfb79;
assign i[5990]= 16'hf91d;
assign i[5991]= 16'hf731;
assign i[5992]= 16'hf5ba;
assign i[5993]= 16'hf4b8;
assign i[5994]= 16'hf42d;
assign i[5995]= 16'hf415;
assign i[5996]= 16'hf46c;
assign i[5997]= 16'hf52c;
assign i[5998]= 16'hf64e;
assign i[5999]= 16'hf7c8;
assign i[6000]= 16'hf990;
assign i[6001]= 16'hfb9c;
assign i[6002]= 16'hfde2;
assign i[6003]= 16'h54;
assign i[6004]= 16'h2eb;
assign i[6005]= 16'h59a;
assign i[6006]= 16'h858;
assign i[6007]= 16'hb1c;
assign i[6008]= 16'hddd;
assign i[6009]= 16'h1093;
assign i[6010]= 16'h1339;
assign i[6011]= 16'h15c8;
assign i[6012]= 16'h183d;
assign i[6013]= 16'h1a93;
assign i[6014]= 16'h1cc7;
assign i[6015]= 16'h1ed8;
assign i[6016]= 16'h20c2;
assign i[6017]= 16'h2286;
assign i[6018]= 16'h2421;
assign i[6019]= 16'h2592;
assign i[6020]= 16'h26d7;
assign i[6021]= 16'h27f0;
assign i[6022]= 16'h28da;
assign i[6023]= 16'h2994;
assign i[6024]= 16'h2a1b;
assign i[6025]= 16'h2a6c;
assign i[6026]= 16'h2a84;
assign i[6027]= 16'h2a5f;
assign i[6028]= 16'h29fc;
assign i[6029]= 16'h2955;
assign i[6030]= 16'h2869;
assign i[6031]= 16'h2734;
assign i[6032]= 16'h25b5;
assign i[6033]= 16'h23e9;
assign i[6034]= 16'h21d0;
assign i[6035]= 16'h1f6b;
assign i[6036]= 16'h1cba;
assign i[6037]= 16'h19c2;
assign i[6038]= 16'h1686;
assign i[6039]= 16'h130b;
assign i[6040]= 16'hf59;
assign i[6041]= 16'hb78;
assign i[6042]= 16'h770;
assign i[6043]= 16'h34c;
assign i[6044]= 16'hff19;
assign i[6045]= 16'hfae0;
assign i[6046]= 16'hf6af;
assign i[6047]= 16'hf292;
assign i[6048]= 16'hee96;
assign i[6049]= 16'heac7;
assign i[6050]= 16'he730;
assign i[6051]= 16'he3dd;
assign i[6052]= 16'he0d7;
assign i[6053]= 16'hde27;
assign i[6054]= 16'hdbd4;
assign i[6055]= 16'hd9e4;
assign i[6056]= 16'hd85c;
assign i[6057]= 16'hd73e;
assign i[6058]= 16'hd68b;
assign i[6059]= 16'hd643;
assign i[6060]= 16'hd662;
assign i[6061]= 16'hd6e6;
assign i[6062]= 16'hd7c9;
assign i[6063]= 16'hd905;
assign i[6064]= 16'hda91;
assign i[6065]= 16'hdc66;
assign i[6066]= 16'hde78;
assign i[6067]= 16'he0bd;
assign i[6068]= 16'he32a;
assign i[6069]= 16'he5b2;
assign i[6070]= 16'he84a;
assign i[6071]= 16'heae4;
assign i[6072]= 16'hed74;
assign i[6073]= 16'hefed;
assign i[6074]= 16'hf242;
assign i[6075]= 16'hf467;
assign i[6076]= 16'hf650;
assign i[6077]= 16'hf7f3;
assign i[6078]= 16'hf945;
assign i[6079]= 16'hfa3d;
assign i[6080]= 16'hfad4;
assign i[6081]= 16'hfb04;
assign i[6082]= 16'hfac9;
assign i[6083]= 16'hfa22;
assign i[6084]= 16'hf90d;
assign i[6085]= 16'hf78f;
assign i[6086]= 16'hf5ad;
assign i[6087]= 16'hf36d;
assign i[6088]= 16'hf0dc;
assign i[6089]= 16'hee07;
assign i[6090]= 16'heafc;
assign i[6091]= 16'he7ce;
assign i[6092]= 16'he491;
assign i[6093]= 16'he15a;
assign i[6094]= 16'hde3f;
assign i[6095]= 16'hdb59;
assign i[6096]= 16'hd8be;
assign i[6097]= 16'hd686;
assign i[6098]= 16'hd4c4;
assign i[6099]= 16'hd38e;
assign i[6100]= 16'hd2f3;
assign i[6101]= 16'hd303;
assign i[6102]= 16'hd3c6;
assign i[6103]= 16'hd544;
assign i[6104]= 16'hd77d;
assign i[6105]= 16'hda6e;
assign i[6106]= 16'hde10;
assign i[6107]= 16'he255;
assign i[6108]= 16'he72b;
assign i[6109]= 16'hec7e;
assign i[6110]= 16'hf232;
assign i[6111]= 16'hf82a;
assign i[6112]= 16'hfe48;
assign i[6113]= 16'h469;
assign i[6114]= 16'ha6d;
assign i[6115]= 16'h1031;
assign i[6116]= 16'h1594;
assign i[6117]= 16'h1a77;
assign i[6118]= 16'h1ebf;
assign i[6119]= 16'h2252;
assign i[6120]= 16'h251e;
assign i[6121]= 16'h2712;
assign i[6122]= 16'h2826;
assign i[6123]= 16'h2855;
assign i[6124]= 16'h27a1;
assign i[6125]= 16'h2611;
assign i[6126]= 16'h23b2;
assign i[6127]= 16'h2094;
assign i[6128]= 16'h1ccc;
assign i[6129]= 16'h1874;
assign i[6130]= 16'h13a7;
assign i[6131]= 16'he82;
assign i[6132]= 16'h924;
assign i[6133]= 16'h3a9;
assign i[6134]= 16'hfe31;
assign i[6135]= 16'hf8d4;
assign i[6136]= 16'hf3ad;
assign i[6137]= 16'heed0;
assign i[6138]= 16'hea50;
assign i[6139]= 16'he63c;
assign i[6140]= 16'he29c;
assign i[6141]= 16'hdf77;
assign i[6142]= 16'hdcd0;
assign i[6143]= 16'hdaa3;
assign i[6144]= 16'hd8ee;
assign i[6145]= 16'hd7a7;
assign i[6146]= 16'hd6c4;
assign i[6147]= 16'hd63c;
assign i[6148]= 16'hd601;
assign i[6149]= 16'hd607;
assign i[6150]= 16'hd643;
assign i[6151]= 16'hd6a9;
assign i[6152]= 16'hd730;
assign i[6153]= 16'hd7d0;
assign i[6154]= 16'hd885;
assign i[6155]= 16'hd949;
assign i[6156]= 16'hda1d;
assign i[6157]= 16'hdb01;
assign i[6158]= 16'hdbf9;
assign i[6159]= 16'hdd07;
assign i[6160]= 16'hde31;
assign i[6161]= 16'hdf7d;
assign i[6162]= 16'he0f1;
assign i[6163]= 16'he291;
assign i[6164]= 16'he463;
assign i[6165]= 16'he669;
assign i[6166]= 16'he8a4;
assign i[6167]= 16'heb13;
assign i[6168]= 16'hedb2;
assign i[6169]= 16'hf07c;
assign i[6170]= 16'hf369;
assign i[6171]= 16'hf66d;
assign i[6172]= 16'hf97d;
assign i[6173]= 16'hfc8a;
assign i[6174]= 16'hff86;
assign i[6175]= 16'h25f;
assign i[6176]= 16'h507;
assign i[6177]= 16'h76f;
assign i[6178]= 16'h988;
assign i[6179]= 16'hb45;
assign i[6180]= 16'hc9c;
assign i[6181]= 16'hd86;
assign i[6182]= 16'hdfd;
assign i[6183]= 16'he01;
assign i[6184]= 16'hd93;
assign i[6185]= 16'hcb8;
assign i[6186]= 16'hb79;
assign i[6187]= 16'h9e1;
assign i[6188]= 16'h7ff;
assign i[6189]= 16'h5e2;
assign i[6190]= 16'h39c;
assign i[6191]= 16'h141;
assign i[6192]= 16'hfee5;
assign i[6193]= 16'hfc99;
assign i[6194]= 16'hfa71;
assign i[6195]= 16'hf87d;
assign i[6196]= 16'hf6cc;
assign i[6197]= 16'hf56d;
assign i[6198]= 16'hf467;
assign i[6199]= 16'hf3c3;
assign i[6200]= 16'hf384;
assign i[6201]= 16'hf3ab;
assign i[6202]= 16'hf434;
assign i[6203]= 16'hf51c;
assign i[6204]= 16'hf659;
assign i[6205]= 16'hf7e0;
assign i[6206]= 16'hf9a6;
assign i[6207]= 16'hfb9d;
assign i[6208]= 16'hfdb6;
assign i[6209]= 16'hffe2;
assign i[6210]= 16'h211;
assign i[6211]= 16'h438;
assign i[6212]= 16'h647;
assign i[6213]= 16'h835;
assign i[6214]= 16'h9f7;
assign i[6215]= 16'hb85;
assign i[6216]= 16'hcdb;
assign i[6217]= 16'hdf7;
assign i[6218]= 16'hed7;
assign i[6219]= 16'hf7e;
assign i[6220]= 16'hfef;
assign i[6221]= 16'h1030;
assign i[6222]= 16'h104a;
assign i[6223]= 16'h1044;
assign i[6224]= 16'h1028;
assign i[6225]= 16'h1000;
assign i[6226]= 16'hfd7;
assign i[6227]= 16'hfb7;
assign i[6228]= 16'hfa8;
assign i[6229]= 16'hfb4;
assign i[6230]= 16'hfe3;
assign i[6231]= 16'h1039;
assign i[6232]= 16'h10bd;
assign i[6233]= 16'h1171;
assign i[6234]= 16'h1256;
assign i[6235]= 16'h136d;
assign i[6236]= 16'h14b4;
assign i[6237]= 16'h1627;
assign i[6238]= 16'h17c1;
assign i[6239]= 16'h197e;
assign i[6240]= 16'h1b54;
assign i[6241]= 16'h1d3d;
assign i[6242]= 16'h1f30;
assign i[6243]= 16'h2122;
assign i[6244]= 16'h230b;
assign i[6245]= 16'h24e0;
assign i[6246]= 16'h2696;
assign i[6247]= 16'h2824;
assign i[6248]= 16'h2980;
assign i[6249]= 16'h2aa0;
assign i[6250]= 16'h2b7b;
assign i[6251]= 16'h2c08;
assign i[6252]= 16'h2c40;
assign i[6253]= 16'h2c1b;
assign i[6254]= 16'h2b95;
assign i[6255]= 16'h2aa7;
assign i[6256]= 16'h294f;
assign i[6257]= 16'h278a;
assign i[6258]= 16'h2558;
assign i[6259]= 16'h22b9;
assign i[6260]= 16'h1fb2;
assign i[6261]= 16'h1c46;
assign i[6262]= 16'h187c;
assign i[6263]= 16'h145e;
assign i[6264]= 16'hff5;
assign i[6265]= 16'hb4f;
assign i[6266]= 16'h67a;
assign i[6267]= 16'h188;
assign i[6268]= 16'hfc8a;
assign i[6269]= 16'hf792;
assign i[6270]= 16'hf2b5;
assign i[6271]= 16'hee09;
assign i[6272]= 16'he9a1;
assign i[6273]= 16'he592;
assign i[6274]= 16'he1ef;
assign i[6275]= 16'hdecb;
assign i[6276]= 16'hdc35;
assign i[6277]= 16'hda3c;
assign i[6278]= 16'hd8e8;
assign i[6279]= 16'hd842;
assign i[6280]= 16'hd84c;
assign i[6281]= 16'hd906;
assign i[6282]= 16'hda6a;
assign i[6283]= 16'hdc71;
assign i[6284]= 16'hdf0c;
assign i[6285]= 16'he22b;
assign i[6286]= 16'he5b8;
assign i[6287]= 16'he99c;
assign i[6288]= 16'hedbe;
assign i[6289]= 16'hf200;
assign i[6290]= 16'hf648;
assign i[6291]= 16'hfa76;
assign i[6292]= 16'hfe70;
assign i[6293]= 16'h21a;
assign i[6294]= 16'h55d;
assign i[6295]= 16'h824;
assign i[6296]= 16'ha5e;
assign i[6297]= 16'hbfe;
assign i[6298]= 16'hcfd;
assign i[6299]= 16'hd57;
assign i[6300]= 16'hd11;
assign i[6301]= 16'hc31;
assign i[6302]= 16'hac4;
assign i[6303]= 16'h8db;
assign i[6304]= 16'h68c;
assign i[6305]= 16'h3ee;
assign i[6306]= 16'h11b;
assign i[6307]= 16'hfe2f;
assign i[6308]= 16'hfb43;
assign i[6309]= 16'hf871;
assign i[6310]= 16'hf5d3;
assign i[6311]= 16'hf37d;
assign i[6312]= 16'hf181;
assign i[6313]= 16'hefea;
assign i[6314]= 16'heec2;
assign i[6315]= 16'hee09;
assign i[6316]= 16'hedbe;
assign i[6317]= 16'hedd8;
assign i[6318]= 16'hee4a;
assign i[6319]= 16'hef02;
assign i[6320]= 16'hefea;
assign i[6321]= 16'hf0ec;
assign i[6322]= 16'hf1ee;
assign i[6323]= 16'hf2d6;
assign i[6324]= 16'hf38a;
assign i[6325]= 16'hf3f4;
assign i[6326]= 16'hf400;
assign i[6327]= 16'hf39f;
assign i[6328]= 16'hf2c4;
assign i[6329]= 16'hf16d;
assign i[6330]= 16'hef99;
assign i[6331]= 16'hed51;
assign i[6332]= 16'heaa1;
assign i[6333]= 16'he79f;
assign i[6334]= 16'he463;
assign i[6335]= 16'he10a;
assign i[6336]= 16'hddb5;
assign i[6337]= 16'hda87;
assign i[6338]= 16'hd7a3;
assign i[6339]= 16'hd52c;
assign i[6340]= 16'hd340;
assign i[6341]= 16'hd1fd;
assign i[6342]= 16'hd179;
assign i[6343]= 16'hd1c4;
assign i[6344]= 16'hd2e8;
assign i[6345]= 16'hd4e5;
assign i[6346]= 16'hd7b4;
assign i[6347]= 16'hdb46;
assign i[6348]= 16'hdf82;
assign i[6349]= 16'he44a;
assign i[6350]= 16'he978;
assign i[6351]= 16'heee0;
assign i[6352]= 16'hf456;
assign i[6353]= 16'hf9a8;
assign i[6354]= 16'hfea7;
assign i[6355]= 16'h322;
assign i[6356]= 16'h6f1;
assign i[6357]= 16'h9ef;
assign i[6358]= 16'hbfc;
assign i[6359]= 16'hd04;
assign i[6360]= 16'hcf9;
assign i[6361]= 16'hbdc;
assign i[6362]= 16'h9b3;
assign i[6363]= 16'h693;
assign i[6364]= 16'h298;
assign i[6365]= 16'hfdea;
assign i[6366]= 16'hf8b4;
assign i[6367]= 16'hf32c;
assign i[6368]= 16'hed8b;
assign i[6369]= 16'he80a;
assign i[6370]= 16'he2e4;
assign i[6371]= 16'hde51;
assign i[6372]= 16'hda85;
assign i[6373]= 16'hd7ad;
assign i[6374]= 16'hd5ec;
assign i[6375]= 16'hd55f;
assign i[6376]= 16'hd614;
assign i[6377]= 16'hd80e;
assign i[6378]= 16'hdb45;
assign i[6379]= 16'hdfa5;
assign i[6380]= 16'he50c;
assign i[6381]= 16'heb50;
assign i[6382]= 16'hf23e;
assign i[6383]= 16'hf99a;
assign i[6384]= 16'h125;
assign i[6385]= 16'h89e;
assign i[6386]= 16'hfc2;
assign i[6387]= 16'h1650;
assign i[6388]= 16'h1c0f;
assign i[6389]= 16'h20c9;
assign i[6390]= 16'h2454;
assign i[6391]= 16'h268f;
assign i[6392]= 16'h2766;
assign i[6393]= 16'h26d1;
assign i[6394]= 16'h24d6;
assign i[6395]= 16'h2186;
assign i[6396]= 16'h1d02;
assign i[6397]= 16'h1773;
assign i[6398]= 16'h110d;
assign i[6399]= 16'ha0b;
assign i[6400]= 16'h2b0;
assign i[6401]= 16'hfb3f;
assign i[6402]= 16'hf3fd;
assign i[6403]= 16'hed2e;
assign i[6404]= 16'he711;
assign i[6405]= 16'he1df;
assign i[6406]= 16'hddc6;
assign i[6407]= 16'hdaed;
assign i[6408]= 16'hd96e;
assign i[6409]= 16'hd954;
assign i[6410]= 16'hdaa1;
assign i[6411]= 16'hdd47;
assign i[6412]= 16'he12d;
assign i[6413]= 16'he62f;
assign i[6414]= 16'hec1d;
assign i[6415]= 16'hf2c0;
assign i[6416]= 16'hf9db;
assign i[6417]= 16'h12c;
assign i[6418]= 16'h871;
assign i[6419]= 16'hf69;
assign i[6420]= 16'h15d3;
assign i[6421]= 16'h1b77;
assign i[6422]= 16'h2022;
assign i[6423]= 16'h23ac;
assign i[6424]= 16'h25f5;
assign i[6425]= 16'h26ea;
assign i[6426]= 16'h2684;
assign i[6427]= 16'h24c8;
assign i[6428]= 16'h21c4;
assign i[6429]= 16'h1d95;
assign i[6430]= 16'h185f;
assign i[6431]= 16'h124f;
assign i[6432]= 16'hb99;
assign i[6433]= 16'h475;
assign i[6434]= 16'hfd1f;
assign i[6435]= 16'hf5d1;
assign i[6436]= 16'heec7;
assign i[6437]= 16'he836;
assign i[6438]= 16'he251;
assign i[6439]= 16'hdd42;
assign i[6440]= 16'hd92e;
assign i[6441]= 16'hd62f;
assign i[6442]= 16'hd455;
assign i[6443]= 16'hd3a7;
assign i[6444]= 16'hd425;
assign i[6445]= 16'hd5c1;
assign i[6446]= 16'hd869;
assign i[6447]= 16'hdc01;
assign i[6448]= 16'he069;
assign i[6449]= 16'he57a;
assign i[6450]= 16'heb0c;
assign i[6451]= 16'hf0f5;
assign i[6452]= 16'hf709;
assign i[6453]= 16'hfd21;
assign i[6454]= 16'h315;
assign i[6455]= 16'h8c6;
assign i[6456]= 16'he16;
assign i[6457]= 16'h12ed;
assign i[6458]= 16'h173c;
assign i[6459]= 16'h1af8;
assign i[6460]= 16'h1e1d;
assign i[6461]= 16'h20af;
assign i[6462]= 16'h22b5;
assign i[6463]= 16'h243c;
assign i[6464]= 16'h2555;
assign i[6465]= 16'h2615;
assign i[6466]= 16'h2690;
assign i[6467]= 16'h26dd;
assign i[6468]= 16'h2712;
assign i[6469]= 16'h2743;
assign i[6470]= 16'h2782;
assign i[6471]= 16'h27dc;
assign i[6472]= 16'h285e;
assign i[6473]= 16'h290c;
assign i[6474]= 16'h29e9;
assign i[6475]= 16'h2af2;
assign i[6476]= 16'h2c1f;
assign i[6477]= 16'h2d66;
assign i[6478]= 16'h2eb8;
assign i[6479]= 16'h3004;
assign i[6480]= 16'h3138;
assign i[6481]= 16'h3241;
assign i[6482]= 16'h330d;
assign i[6483]= 16'h3388;
assign i[6484]= 16'h33a6;
assign i[6485]= 16'h3359;
assign i[6486]= 16'h3299;
assign i[6487]= 16'h3163;
assign i[6488]= 16'h2fb7;
assign i[6489]= 16'h2d9c;
assign i[6490]= 16'h2b1c;
assign i[6491]= 16'h2848;
assign i[6492]= 16'h2532;
assign i[6493]= 16'h21f1;
assign i[6494]= 16'h1ea1;
assign i[6495]= 16'h1b5c;
assign i[6496]= 16'h183e;
assign i[6497]= 16'h1564;
assign i[6498]= 16'h12e7;
assign i[6499]= 16'h10e0;
assign i[6500]= 16'hf60;
assign i[6501]= 16'he79;
assign i[6502]= 16'he33;
assign i[6503]= 16'he93;
assign i[6504]= 16'hf95;
assign i[6505]= 16'h1130;
assign i[6506]= 16'h1357;
assign i[6507]= 16'h15f3;
assign i[6508]= 16'h18ec;
assign i[6509]= 16'h1c21;
assign i[6510]= 16'h1f71;
assign i[6511]= 16'h22b8;
assign i[6512]= 16'h25d2;
assign i[6513]= 16'h2898;
assign i[6514]= 16'h2ae8;
assign i[6515]= 16'h2ca3;
assign i[6516]= 16'h2dac;
assign i[6517]= 16'h2dec;
assign i[6518]= 16'h2d54;
assign i[6519]= 16'h2bd9;
assign i[6520]= 16'h297b;
assign i[6521]= 16'h263e;
assign i[6522]= 16'h222f;
assign i[6523]= 16'h1d62;
assign i[6524]= 16'h17f2;
assign i[6525]= 16'h1200;
assign i[6526]= 16'hbb1;
assign i[6527]= 16'h52d;
assign i[6528]= 16'hfea1;
assign i[6529]= 16'hf836;
assign i[6530]= 16'hf21b;
assign i[6531]= 16'hec77;
assign i[6532]= 16'he773;
assign i[6533]= 16'he330;
assign i[6534]= 16'hdfcc;
assign i[6535]= 16'hdd5e;
assign i[6536]= 16'hdbf5;
assign i[6537]= 16'hdb9c;
assign i[6538]= 16'hdc52;
assign i[6539]= 16'hde13;
assign i[6540]= 16'he0d2;
assign i[6541]= 16'he47c;
assign i[6542]= 16'he8f8;
assign i[6543]= 16'hee27;
assign i[6544]= 16'hf3ea;
assign i[6545]= 16'hfa1a;
assign i[6546]= 16'h90;
assign i[6547]= 16'h728;
assign i[6548]= 16'hdb9;
assign i[6549]= 16'h141e;
assign i[6550]= 16'h1a34;
assign i[6551]= 16'h1fd9;
assign i[6552]= 16'h24f2;
assign i[6553]= 16'h2966;
assign i[6554]= 16'h2d20;
assign i[6555]= 16'h3010;
assign i[6556]= 16'h322c;
assign i[6557]= 16'h336d;
assign i[6558]= 16'h33d1;
assign i[6559]= 16'h335b;
assign i[6560]= 16'h320f;
assign i[6561]= 16'h2ff7;
assign i[6562]= 16'h2d21;
assign i[6563]= 16'h299b;
assign i[6564]= 16'h2577;
assign i[6565]= 16'h20c7;
assign i[6566]= 16'h1ba3;
assign i[6567]= 16'h1620;
assign i[6568]= 16'h1055;
assign i[6569]= 16'ha5b;
assign i[6570]= 16'h44b;
assign i[6571]= 16'hfe40;
assign i[6572]= 16'hf851;
assign i[6573]= 16'hf298;
assign i[6574]= 16'hed2d;
assign i[6575]= 16'he82a;
assign i[6576]= 16'he3a4;
assign i[6577]= 16'hdfb2;
assign i[6578]= 16'hdc66;
assign i[6579]= 16'hd9d2;
assign i[6580]= 16'hd804;
assign i[6581]= 16'hd708;
assign i[6582]= 16'hd6e3;
assign i[6583]= 16'hd79b;
assign i[6584]= 16'hd92c;
assign i[6585]= 16'hdb93;
assign i[6586]= 16'hdec3;
assign i[6587]= 16'he2ae;
assign i[6588]= 16'he741;
assign i[6589]= 16'hec63;
assign i[6590]= 16'hf1f8;
assign i[6591]= 16'hf7e3;
assign i[6592]= 16'hfe02;
assign i[6593]= 16'h430;
assign i[6594]= 16'ha4e;
assign i[6595]= 16'h1038;
assign i[6596]= 16'h15cb;
assign i[6597]= 16'h1aeb;
assign i[6598]= 16'h1f7a;
assign i[6599]= 16'h2363;
assign i[6600]= 16'h2693;
assign i[6601]= 16'h2900;
assign i[6602]= 16'h2aa1;
assign i[6603]= 16'h2b79;
assign i[6604]= 16'h2b8d;
assign i[6605]= 16'h2ae9;
assign i[6606]= 16'h29a0;
assign i[6607]= 16'h27c7;
assign i[6608]= 16'h2578;
assign i[6609]= 16'h22d2;
assign i[6610]= 16'h1ff2;
assign i[6611]= 16'h1cf7;
assign i[6612]= 16'h19ff;
assign i[6613]= 16'h1728;
assign i[6614]= 16'h148a;
assign i[6615]= 16'h123b;
assign i[6616]= 16'h104b;
assign i[6617]= 16'hec6;
assign i[6618]= 16'hdb0;
assign i[6619]= 16'hd09;
assign i[6620]= 16'hccc;
assign i[6621]= 16'hcec;
assign i[6622]= 16'hd59;
assign i[6623]= 16'hdff;
assign i[6624]= 16'hec6;
assign i[6625]= 16'hf96;
assign i[6626]= 16'h1054;
assign i[6627]= 16'h10e5;
assign i[6628]= 16'h1132;
assign i[6629]= 16'h1125;
assign i[6630]= 16'h10ab;
assign i[6631]= 16'hfb7;
assign i[6632]= 16'he3f;
assign i[6633]= 16'hc40;
assign i[6634]= 16'h9bb;
assign i[6635]= 16'h6b8;
assign i[6636]= 16'h344;
assign i[6637]= 16'hff6f;
assign i[6638]= 16'hfb4e;
assign i[6639]= 16'hf6fb;
assign i[6640]= 16'hf28f;
assign i[6641]= 16'hee27;
assign i[6642]= 16'he9e0;
assign i[6643]= 16'he5d6;
assign i[6644]= 16'he223;
assign i[6645]= 16'hdedf;
assign i[6646]= 16'hdc20;
assign i[6647]= 16'hd9f6;
assign i[6648]= 16'hd870;
assign i[6649]= 16'hd796;
assign i[6650]= 16'hd76e;
assign i[6651]= 16'hd7f8;
assign i[6652]= 16'hd931;
assign i[6653]= 16'hdb11;
assign i[6654]= 16'hdd8f;
assign i[6655]= 16'he09e;
assign i[6656]= 16'he430;
assign i[6657]= 16'he833;
assign i[6658]= 16'hec96;
assign i[6659]= 16'hf148;
assign i[6660]= 16'hf636;
assign i[6661]= 16'hfb4d;
assign i[6662]= 16'h7b;
assign i[6663]= 16'h5b1;
assign i[6664]= 16'hadd;
assign i[6665]= 16'hfee;
assign i[6666]= 16'h14d5;
assign i[6667]= 16'h1983;
assign i[6668]= 16'h1de9;
assign i[6669]= 16'h21f9;
assign i[6670]= 16'h25a4;
assign i[6671]= 16'h28de;
assign i[6672]= 16'h2b99;
assign i[6673]= 16'h2dca;
assign i[6674]= 16'h2f64;
assign i[6675]= 16'h3060;
assign i[6676]= 16'h30b4;
assign i[6677]= 16'h305d;
assign i[6678]= 16'h2f58;
assign i[6679]= 16'h2da7;
assign i[6680]= 16'h2b4d;
assign i[6681]= 16'h2855;
assign i[6682]= 16'h24cc;
assign i[6683]= 16'h20c5;
assign i[6684]= 16'h1c55;
assign i[6685]= 16'h1799;
assign i[6686]= 16'h12ad;
assign i[6687]= 16'hdb3;
assign i[6688]= 16'h8cf;
assign i[6689]= 16'h426;
assign i[6690]= 16'hffdc;
assign i[6691]= 16'hfc14;
assign i[6692]= 16'hf8ee;
assign i[6693]= 16'hf686;
assign i[6694]= 16'hf4f5;
assign i[6695]= 16'hf44b;
assign i[6696]= 16'hf492;
assign i[6697]= 16'hf5ca;
assign i[6698]= 16'hf7ed;
assign i[6699]= 16'hfaeb;
assign i[6700]= 16'hfeac;
assign i[6701]= 16'h30e;
assign i[6702]= 16'h7ec;
assign i[6703]= 16'hd18;
assign i[6704]= 16'h1260;
assign i[6705]= 16'h1791;
assign i[6706]= 16'h1c73;
assign i[6707]= 16'h20d4;
assign i[6708]= 16'h2483;
assign i[6709]= 16'h2754;
assign i[6710]= 16'h2922;
assign i[6711]= 16'h29d0;
assign i[6712]= 16'h294d;
assign i[6713]= 16'h2792;
assign i[6714]= 16'h24a2;
assign i[6715]= 16'h208d;
assign i[6716]= 16'h1b6e;
assign i[6717]= 16'h156c;
assign i[6718]= 16'heb6;
assign i[6719]= 16'h782;
assign i[6720]= 16'hd;
assign i[6721]= 16'hf899;
assign i[6722]= 16'hf166;
assign i[6723]= 16'heab5;
assign i[6724]= 16'he4c4;
assign i[6725]= 16'hdfca;
assign i[6726]= 16'hdbf5;
assign i[6727]= 16'hd96a;
assign i[6728]= 16'hd842;
assign i[6729]= 16'hd889;
assign i[6730]= 16'hda3f;
assign i[6731]= 16'hdd55;
assign i[6732]= 16'he1af;
assign i[6733]= 16'he725;
assign i[6734]= 16'hed86;
assign i[6735]= 16'hf497;
assign i[6736]= 16'hfc14;
assign i[6737]= 16'h3b8;
assign i[6738]= 16'hb3b;
assign i[6739]= 16'h1258;
assign i[6740]= 16'h18ca;
assign i[6741]= 16'h1e55;
assign i[6742]= 16'h22c4;
assign i[6743]= 16'h25ef;
assign i[6744]= 16'h27b7;
assign i[6745]= 16'h280c;
assign i[6746]= 16'h26ec;
assign i[6747]= 16'h2460;
assign i[6748]= 16'h2081;
assign i[6749]= 16'h1b74;
assign i[6750]= 16'h1568;
assign i[6751]= 16'he95;
assign i[6752]= 16'h739;
assign i[6753]= 16'hff99;
assign i[6754]= 16'hf7f8;
assign i[6755]= 16'hf09a;
assign i[6756]= 16'he9c0;
assign i[6757]= 16'he3a4;
assign i[6758]= 16'hde78;
assign i[6759]= 16'hda64;
assign i[6760]= 16'hd787;
assign i[6761]= 16'hd5f0;
assign i[6762]= 16'hd5a5;
assign i[6763]= 16'hd69c;
assign i[6764]= 16'hd8c2;
assign i[6765]= 16'hdbf6;
assign i[6766]= 16'he010;
assign i[6767]= 16'he4df;
assign i[6768]= 16'hea2b;
assign i[6769]= 16'hefb9;
assign i[6770]= 16'hf54e;
assign i[6771]= 16'hfaaf;
assign i[6772]= 16'hffa3;
assign i[6773]= 16'h3f9;
assign i[6774]= 16'h786;
assign i[6775]= 16'ha27;
assign i[6776]= 16'hbc4;
assign i[6777]= 16'hc4f;
assign i[6778]= 16'hbc7;
assign i[6779]= 16'ha31;
assign i[6780]= 16'h7a2;
assign i[6781]= 16'h436;
assign i[6782]= 16'hf;
assign i[6783]= 16'hfb5a;
assign i[6784]= 16'hf645;
assign i[6785]= 16'hf102;
assign i[6786]= 16'hebc6;
assign i[6787]= 16'he6c1;
assign i[6788]= 16'he225;
assign i[6789]= 16'hde1b;
assign i[6790]= 16'hdac8;
assign i[6791]= 16'hd84a;
assign i[6792]= 16'hd6b5;
assign i[6793]= 16'hd615;
assign i[6794]= 16'hd66f;
assign i[6795]= 16'hd7bb;
assign i[6796]= 16'hd9ec;
assign i[6797]= 16'hdcec;
assign i[6798]= 16'he09e;
assign i[6799]= 16'he4e0;
assign i[6800]= 16'he98b;
assign i[6801]= 16'hee77;
assign i[6802]= 16'hf37b;
assign i[6803]= 16'hf86c;
assign i[6804]= 16'hfd24;
assign i[6805]= 16'h17e;
assign i[6806]= 16'h55c;
assign i[6807]= 16'h8a4;
assign i[6808]= 16'hb42;
assign i[6809]= 16'hd28;
assign i[6810]= 16'he51;
assign i[6811]= 16'hebd;
assign i[6812]= 16'he72;
assign i[6813]= 16'hd7f;
assign i[6814]= 16'hbf4;
assign i[6815]= 16'h9ea;
assign i[6816]= 16'h77a;
assign i[6817]= 16'h4c0;
assign i[6818]= 16'h1db;
assign i[6819]= 16'hfee9;
assign i[6820]= 16'hfc06;
assign i[6821]= 16'hf94f;
assign i[6822]= 16'hf6dc;
assign i[6823]= 16'hf4c2;
assign i[6824]= 16'hf315;
assign i[6825]= 16'hf1e0;
assign i[6826]= 16'hf12e;
assign i[6827]= 16'hf102;
assign i[6828]= 16'hf15e;
assign i[6829]= 16'hf23c;
assign i[6830]= 16'hf396;
assign i[6831]= 16'hf561;
assign i[6832]= 16'hf78e;
assign i[6833]= 16'hfa0f;
assign i[6834]= 16'hfcd2;
assign i[6835]= 16'hffc7;
assign i[6836]= 16'h2d9;
assign i[6837]= 16'h5fb;
assign i[6838]= 16'h91c;
assign i[6839]= 16'hc2d;
assign i[6840]= 16'hf22;
assign i[6841]= 16'h11f1;
assign i[6842]= 16'h1494;
assign i[6843]= 16'h1704;
assign i[6844]= 16'h1940;
assign i[6845]= 16'h1b48;
assign i[6846]= 16'h1d1d;
assign i[6847]= 16'h1ec5;
assign i[6848]= 16'h2044;
assign i[6849]= 16'h21a1;
assign i[6850]= 16'h22e4;
assign i[6851]= 16'h2413;
assign i[6852]= 16'h2536;
assign i[6853]= 16'h2654;
assign i[6854]= 16'h2772;
assign i[6855]= 16'h2893;
assign i[6856]= 16'h29bb;
assign i[6857]= 16'h2ae9;
assign i[6858]= 16'h2c1c;
assign i[6859]= 16'h2d50;
assign i[6860]= 16'h2e81;
assign i[6861]= 16'h2fa5;
assign i[6862]= 16'h30b5;
assign i[6863]= 16'h31a7;
assign i[6864]= 16'h326f;
assign i[6865]= 16'h3304;
assign i[6866]= 16'h3359;
assign i[6867]= 16'h3366;
assign i[6868]= 16'h3322;
assign i[6869]= 16'h3287;
assign i[6870]= 16'h318f;
assign i[6871]= 16'h3039;
assign i[6872]= 16'h2e88;
assign i[6873]= 16'h2c7f;
assign i[6874]= 16'h2a27;
assign i[6875]= 16'h278c;
assign i[6876]= 16'h24bc;
assign i[6877]= 16'h21c9;
assign i[6878]= 16'h1ec7;
assign i[6879]= 16'h1bcb;
assign i[6880]= 16'h18ed;
assign i[6881]= 16'h1644;
assign i[6882]= 16'h13e7;
assign i[6883]= 16'h11eb;
assign i[6884]= 16'h1063;
assign i[6885]= 16'hf5e;
assign i[6886]= 16'hee9;
assign i[6887]= 16'hf0b;
assign i[6888]= 16'hfc6;
assign i[6889]= 16'h1115;
assign i[6890]= 16'h12ef;
assign i[6891]= 16'h1545;
assign i[6892]= 16'h1803;
assign i[6893]= 16'h1b0d;
assign i[6894]= 16'h1e46;
assign i[6895]= 16'h218c;
assign i[6896]= 16'h24ba;
assign i[6897]= 16'h27ac;
assign i[6898]= 16'h2a3c;
assign i[6899]= 16'h2c47;
assign i[6900]= 16'h2dac;
assign i[6901]= 16'h2e4e;
assign i[6902]= 16'h2e17;
assign i[6903]= 16'h2cf6;
assign i[6904]= 16'h2ae3;
assign i[6905]= 16'h27dd;
assign i[6906]= 16'h23ec;
assign i[6907]= 16'h1f1f;
assign i[6908]= 16'h1991;
assign i[6909]= 16'h1360;
assign i[6910]= 16'hcb4;
assign i[6911]= 16'h5b8;
assign i[6912]= 16'hfe9e;
assign i[6913]= 16'hf797;
assign i[6914]= 16'hf0d6;
assign i[6915]= 16'hea8e;
assign i[6916]= 16'he4ed;
assign i[6917]= 16'he01d;
assign i[6918]= 16'hdc41;
assign i[6919]= 16'hd975;
assign i[6920]= 16'hd7ca;
assign i[6921]= 16'hd74a;
assign i[6922]= 16'hd7f1;
assign i[6923]= 16'hd9b2;
assign i[6924]= 16'hdc78;
assign i[6925]= 16'he021;
assign i[6926]= 16'he485;
assign i[6927]= 16'he974;
assign i[6928]= 16'heeb9;
assign i[6929]= 16'hf41d;
assign i[6930]= 16'hf967;
assign i[6931]= 16'hfe5f;
assign i[6932]= 16'h2d0;
assign i[6933]= 16'h68c;
assign i[6934]= 16'h96b;
assign i[6935]= 16'hb4e;
assign i[6936]= 16'hc21;
assign i[6937]= 16'hbd9;
assign i[6938]= 16'ha79;
assign i[6939]= 16'h80d;
assign i[6940]= 16'h4ae;
assign i[6941]= 16'h7e;
assign i[6942]= 16'hfbab;
assign i[6943]= 16'hf664;
assign i[6944]= 16'hf0e2;
assign i[6945]= 16'heb61;
assign i[6946]= 16'he61c;
assign i[6947]= 16'he14d;
assign i[6948]= 16'hdd2b;
assign i[6949]= 16'hd9e5;
assign i[6950]= 16'hd7a5;
assign i[6951]= 16'hd688;
assign i[6952]= 16'hd6a3;
assign i[6953]= 16'hd7fd;
assign i[6954]= 16'hda93;
assign i[6955]= 16'hde55;
assign i[6956]= 16'he327;
assign i[6957]= 16'he8e4;
assign i[6958]= 16'hef5c;
assign i[6959]= 16'hf659;
assign i[6960]= 16'hfda1;
assign i[6961]= 16'h4f3;
assign i[6962]= 16'hc11;
assign i[6963]= 16'h12bf;
assign i[6964]= 16'h18c1;
assign i[6965]= 16'h1de4;
assign i[6966]= 16'h21fc;
assign i[6967]= 16'h24e7;
assign i[6968]= 16'h268b;
assign i[6969]= 16'h26dd;
assign i[6970]= 16'h25dc;
assign i[6971]= 16'h2391;
assign i[6972]= 16'h2012;
assign i[6973]= 16'h1b7f;
assign i[6974]= 16'h1600;
assign i[6975]= 16'hfc5;
assign i[6976]= 16'h902;
assign i[6977]= 16'h1f1;
assign i[6978]= 16'hfacb;
assign i[6979]= 16'hf3c8;
assign i[6980]= 16'hed1f;
assign i[6981]= 16'he704;
assign i[6982]= 16'he1a2;
assign i[6983]= 16'hdd1e;
assign i[6984]= 16'hd995;
assign i[6985]= 16'hd71c;
assign i[6986]= 16'hd5bc;
assign i[6987]= 16'hd577;
assign i[6988]= 16'hd647;
assign i[6989]= 16'hd81a;
assign i[6990]= 16'hdadc;
assign i[6991]= 16'hde6e;
assign i[6992]= 16'he2ae;
assign i[6993]= 16'he779;
assign i[6994]= 16'heca6;
assign i[6995]= 16'hf20e;
assign i[6996]= 16'hf78a;
assign i[6997]= 16'hfcf4;
assign i[6998]= 16'h22a;
assign i[6999]= 16'h710;
assign i[7000]= 16'hb8b;
assign i[7001]= 16'hf86;
assign i[7002]= 16'h12f3;
assign i[7003]= 16'h15c8;
assign i[7004]= 16'h17ff;
assign i[7005]= 16'h1998;
assign i[7006]= 16'h1a98;
assign i[7007]= 16'h1b06;
assign i[7008]= 16'h1aed;
assign i[7009]= 16'h1a5a;
assign i[7010]= 16'h195b;
assign i[7011]= 16'h17ff;
assign i[7012]= 16'h1657;
assign i[7013]= 16'h1472;
assign i[7014]= 16'h125e;
assign i[7015]= 16'h1029;
assign i[7016]= 16'hddf;
assign i[7017]= 16'hb8c;
assign i[7018]= 16'h939;
assign i[7019]= 16'h6ee;
assign i[7020]= 16'h4b2;
assign i[7021]= 16'h289;
assign i[7022]= 16'h7a;
assign i[7023]= 16'hfe88;
assign i[7024]= 16'hfcb3;
assign i[7025]= 16'hfb00;
assign i[7026]= 16'hf96f;
assign i[7027]= 16'hf803;
assign i[7028]= 16'hf6bc;
assign i[7029]= 16'hf59a;
assign i[7030]= 16'hf49e;
assign i[7031]= 16'hf3c8;
assign i[7032]= 16'hf317;
assign i[7033]= 16'hf289;
assign i[7034]= 16'hf21d;
assign i[7035]= 16'hf1d0;
assign i[7036]= 16'hf19d;
assign i[7037]= 16'hf183;
assign i[7038]= 16'hf17a;
assign i[7039]= 16'hf180;
assign i[7040]= 16'hf18d;
assign i[7041]= 16'hf19c;
assign i[7042]= 16'hf1a9;
assign i[7043]= 16'hf1ac;
assign i[7044]= 16'hf1a3;
assign i[7045]= 16'hf189;
assign i[7046]= 16'hf15b;
assign i[7047]= 16'hf118;
assign i[7048]= 16'hf0c1;
assign i[7049]= 16'hf056;
assign i[7050]= 16'hefdc;
assign i[7051]= 16'hef57;
assign i[7052]= 16'heecc;
assign i[7053]= 16'hee45;
assign i[7054]= 16'hedca;
assign i[7055]= 16'hed63;
assign i[7056]= 16'hed1c;
assign i[7057]= 16'hecfe;
assign i[7058]= 16'hed12;
assign i[7059]= 16'hed62;
assign i[7060]= 16'hedf6;
assign i[7061]= 16'heed5;
assign i[7062]= 16'hf003;
assign i[7063]= 16'hf183;
assign i[7064]= 16'hf358;
assign i[7065]= 16'hf580;
assign i[7066]= 16'hf7f8;
assign i[7067]= 16'hfabb;
assign i[7068]= 16'hfdc3;
assign i[7069]= 16'h106;
assign i[7070]= 16'h47c;
assign i[7071]= 16'h818;
assign i[7072]= 16'hbcf;
assign i[7073]= 16'hf92;
assign i[7074]= 16'h1356;
assign i[7075]= 16'h170b;
assign i[7076]= 16'h1aa5;
assign i[7077]= 16'h1e15;
assign i[7078]= 16'h2150;
assign i[7079]= 16'h2448;
assign i[7080]= 16'h26f1;
assign i[7081]= 16'h2941;
assign i[7082]= 16'h2b2d;
assign i[7083]= 16'h2cac;
assign i[7084]= 16'h2db5;
assign i[7085]= 16'h2e41;
assign i[7086]= 16'h2e49;
assign i[7087]= 16'h2dc9;
assign i[7088]= 16'h2cbb;
assign i[7089]= 16'h2b1f;
assign i[7090]= 16'h28f4;
assign i[7091]= 16'h263a;
assign i[7092]= 16'h22f5;
assign i[7093]= 16'h1f2c;
assign i[7094]= 16'h1ae8;
assign i[7095]= 16'h1633;
assign i[7096]= 16'h111c;
assign i[7097]= 16'hbb4;
assign i[7098]= 16'h60f;
assign i[7099]= 16'h45;
assign i[7100]= 16'hfa70;
assign i[7101]= 16'hf4a9;
assign i[7102]= 16'hef0e;
assign i[7103]= 16'he9be;
assign i[7104]= 16'he4d7;
assign i[7105]= 16'he075;
assign i[7106]= 16'hdcb6;
assign i[7107]= 16'hd9b4;
assign i[7108]= 16'hd784;
assign i[7109]= 16'hd638;
assign i[7110]= 16'hd5df;
assign i[7111]= 16'hd680;
assign i[7112]= 16'hd81b;
assign i[7113]= 16'hdaac;
assign i[7114]= 16'hde27;
assign i[7115]= 16'he278;
assign i[7116]= 16'he787;
assign i[7117]= 16'hed34;
assign i[7118]= 16'hf35a;
assign i[7119]= 16'hf9d2;
assign i[7120]= 16'h6e;
assign i[7121]= 16'h702;
assign i[7122]= 16'hd61;
assign i[7123]= 16'h135d;
assign i[7124]= 16'h18cc;
assign i[7125]= 16'h1d88;
assign i[7126]= 16'h2170;
assign i[7127]= 16'h246b;
assign i[7128]= 16'h2665;
assign i[7129]= 16'h2755;
assign i[7130]= 16'h2739;
assign i[7131]= 16'h2618;
assign i[7132]= 16'h2401;
assign i[7133]= 16'h210e;
assign i[7134]= 16'h1d5e;
assign i[7135]= 16'h1917;
assign i[7136]= 16'h1464;
assign i[7137]= 16'hf73;
assign i[7138]= 16'ha76;
assign i[7139]= 16'h59c;
assign i[7140]= 16'h116;
assign i[7141]= 16'hfd10;
assign i[7142]= 16'hf9af;
assign i[7143]= 16'hf716;
assign i[7144]= 16'hf55d;
assign i[7145]= 16'hf495;
assign i[7146]= 16'hf4c8;
assign i[7147]= 16'hf5f3;
assign i[7148]= 16'hf80e;
assign i[7149]= 16'hfb03;
assign i[7150]= 16'hfeba;
assign i[7151]= 16'h310;
assign i[7152]= 16'h7de;
assign i[7153]= 16'hcf9;
assign i[7154]= 16'h1234;
assign i[7155]= 16'h1760;
assign i[7156]= 16'h1c51;
assign i[7157]= 16'h20dc;
assign i[7158]= 16'h24dc;
assign i[7159]= 16'h2831;
assign i[7160]= 16'h2ac2;
assign i[7161]= 16'h2c81;
assign i[7162]= 16'h2d63;
assign i[7163]= 16'h2d6b;
assign i[7164]= 16'h2ca2;
assign i[7165]= 16'h2b19;
assign i[7166]= 16'h28ea;
assign i[7167]= 16'h2634;
assign i[7168]= 16'h231b;
assign i[7169]= 16'h1fc7;
assign i[7170]= 16'h1c63;
assign i[7171]= 16'h1916;
assign i[7172]= 16'h160a;
assign i[7173]= 16'h1363;
assign i[7174]= 16'h1140;
assign i[7175]= 16'hfbb;
assign i[7176]= 16'hee6;
assign i[7177]= 16'hecb;
assign i[7178]= 16'hf6c;
assign i[7179]= 16'h10c2;
assign i[7180]= 16'h12bd;
assign i[7181]= 16'h1547;
assign i[7182]= 16'h1841;
assign i[7183]= 16'h1b89;
assign i[7184]= 16'h1ef6;
assign i[7185]= 16'h225f;
assign i[7186]= 16'h2599;
assign i[7187]= 16'h2879;
assign i[7188]= 16'h2ada;
assign i[7189]= 16'h2c98;
assign i[7190]= 16'h2d97;
assign i[7191]= 16'h2dc1;
assign i[7192]= 16'h2d0a;
assign i[7193]= 16'h2b6d;
assign i[7194]= 16'h28f0;
assign i[7195]= 16'h25a1;
assign i[7196]= 16'h2198;
assign i[7197]= 16'h1cf3;
assign i[7198]= 16'h17d9;
assign i[7199]= 16'h1277;
assign i[7200]= 16'hcfb;
assign i[7201]= 16'h798;
assign i[7202]= 16'h27f;
assign i[7203]= 16'hfde2;
assign i[7204]= 16'hf9eb;
assign i[7205]= 16'hf6c3;
assign i[7206]= 16'hf488;
assign i[7207]= 16'hf352;
assign i[7208]= 16'hf32d;
assign i[7209]= 16'hf41e;
assign i[7210]= 16'hf61c;
assign i[7211]= 16'hf915;
assign i[7212]= 16'hfced;
assign i[7213]= 16'h17e;
assign i[7214]= 16'h69c;
assign i[7215]= 16'hc12;
assign i[7216]= 16'h11a9;
assign i[7217]= 16'h1727;
assign i[7218]= 16'h1c51;
assign i[7219]= 16'h20f0;
assign i[7220]= 16'h24cf;
assign i[7221]= 16'h27c1;
assign i[7222]= 16'h29a0;
assign i[7223]= 16'h2a51;
assign i[7224]= 16'h29c3;
assign i[7225]= 16'h27f2;
assign i[7226]= 16'h24e4;
assign i[7227]= 16'h20ac;
assign i[7228]= 16'h1b6a;
assign i[7229]= 16'h1546;
assign i[7230]= 16'he72;
assign i[7231]= 16'h728;
assign i[7232]= 16'hffa7;
assign i[7233]= 16'hf82f;
assign i[7234]= 16'hf102;
assign i[7235]= 16'hea61;
assign i[7236]= 16'he488;
assign i[7237]= 16'hdfab;
assign i[7238]= 16'hdbf7;
assign i[7239]= 16'hd98e;
assign i[7240]= 16'hd886;
assign i[7241]= 16'hd8ea;
assign i[7242]= 16'hdab6;
assign i[7243]= 16'hddda;
assign i[7244]= 16'he239;
assign i[7245]= 16'he7aa;
assign i[7246]= 16'hedfc;
assign i[7247]= 16'hf4f4;
assign i[7248]= 16'hfc51;
assign i[7249]= 16'h3cf;
assign i[7250]= 16'hb2b;
assign i[7251]= 16'h121e;
assign i[7252]= 16'h186a;
assign i[7253]= 16'h1dd4;
assign i[7254]= 16'h222b;
assign i[7255]= 16'h2547;
assign i[7256]= 16'h270c;
assign i[7257]= 16'h276b;
assign i[7258]= 16'h2661;
assign i[7259]= 16'h23f9;
assign i[7260]= 16'h204a;
assign i[7261]= 16'h1b75;
assign i[7262]= 16'h15a6;
assign i[7263]= 16'hf14;
assign i[7264]= 16'h7f7;
assign i[7265]= 16'h90;
assign i[7266]= 16'hf921;
assign i[7267]= 16'hf1e6;
assign i[7268]= 16'heb1d;
assign i[7269]= 16'he4ff;
assign i[7270]= 16'hdfbb;
assign i[7271]= 16'hdb79;
assign i[7272]= 16'hd857;
assign i[7273]= 16'hd665;
assign i[7274]= 16'hd5ad;
assign i[7275]= 16'hd628;
assign i[7276]= 16'hd7c8;
assign i[7277]= 16'hda73;
assign i[7278]= 16'hde07;
assign i[7279]= 16'he25b;
assign i[7280]= 16'he740;
assign i[7281]= 16'hec83;
assign i[7282]= 16'hf1f1;
assign i[7283]= 16'hf756;
assign i[7284]= 16'hfc82;
assign i[7285]= 16'h146;
assign i[7286]= 16'h57e;
assign i[7287]= 16'h909;
assign i[7288]= 16'hbcf;
assign i[7289]= 16'hdc2;
assign i[7290]= 16'hedc;
assign i[7291]= 16'hf1f;
assign i[7292]= 16'he96;
assign i[7293]= 16'hd55;
assign i[7294]= 16'hb74;
assign i[7295]= 16'h913;
assign i[7296]= 16'h653;
assign i[7297]= 16'h35b;
assign i[7298]= 16'h51;
assign i[7299]= 16'hfd5a;
assign i[7300]= 16'hfa9a;
assign i[7301]= 16'hf831;
assign i[7302]= 16'hf63c;
assign i[7303]= 16'hf4d3;
assign i[7304]= 16'hf408;
assign i[7305]= 16'hf3e7;
assign i[7306]= 16'hf475;
assign i[7307]= 16'hf5b4;
assign i[7308]= 16'hf79d;
assign i[7309]= 16'hfa26;
assign i[7310]= 16'hfd41;
assign i[7311]= 16'hda;
assign i[7312]= 16'h4de;
assign i[7313]= 16'h936;
assign i[7314]= 16'hdca;
assign i[7315]= 16'h1282;
assign i[7316]= 16'h1745;
assign i[7317]= 16'h1bff;
assign i[7318]= 16'h209a;
assign i[7319]= 16'h2501;
assign i[7320]= 16'h2926;
assign i[7321]= 16'h2cf7;
assign i[7322]= 16'h3069;
assign i[7323]= 16'h3370;
assign i[7324]= 16'h3603;
assign i[7325]= 16'h381b;
assign i[7326]= 16'h39b1;
assign i[7327]= 16'h3ac0;
assign i[7328]= 16'h3b45;
assign i[7329]= 16'h3b3c;
assign i[7330]= 16'h3aa4;
assign i[7331]= 16'h397b;
assign i[7332]= 16'h37c1;
assign i[7333]= 16'h3578;
assign i[7334]= 16'h32a1;
assign i[7335]= 16'h2f42;
assign i[7336]= 16'h2b5e;
assign i[7337]= 16'h2700;
assign i[7338]= 16'h222f;
assign i[7339]= 16'h1cfa;
assign i[7340]= 16'h176f;
assign i[7341]= 16'h119e;
assign i[7342]= 16'hb9c;
assign i[7343]= 16'h57c;
assign i[7344]= 16'hff56;
assign i[7345]= 16'hf940;
assign i[7346]= 16'hf351;
assign i[7347]= 16'heda0;
assign i[7348]= 16'he844;
assign i[7349]= 16'he34f;
assign i[7350]= 16'hded4;
assign i[7351]= 16'hdadf;
assign i[7352]= 16'hd77c;
assign i[7353]= 16'hd4b0;
assign i[7354]= 16'hd27c;
assign i[7355]= 16'hd0dd;
assign i[7356]= 16'hcfcc;
assign i[7357]= 16'hcf3c;
assign i[7358]= 16'hcf1d;
assign i[7359]= 16'hcf5d;
assign i[7360]= 16'hcfe6;
assign i[7361]= 16'hd0a0;
assign i[7362]= 16'hd174;
assign i[7363]= 16'hd24b;
assign i[7364]= 16'hd30f;
assign i[7365]= 16'hd3ac;
assign i[7366]= 16'hd414;
assign i[7367]= 16'hd439;
assign i[7368]= 16'hd415;
assign i[7369]= 16'hd3a6;
assign i[7370]= 16'hd2ef;
assign i[7371]= 16'hd1f9;
assign i[7372]= 16'hd0d1;
assign i[7373]= 16'hcf8a;
assign i[7374]= 16'hce38;
assign i[7375]= 16'hccf6;
assign i[7376]= 16'hcbdd;
assign i[7377]= 16'hcb08;
assign i[7378]= 16'hca94;
assign i[7379]= 16'hca98;
assign i[7380]= 16'hcb2c;
assign i[7381]= 16'hcc61;
assign i[7382]= 16'hce46;
assign i[7383]= 16'hd0e2;
assign i[7384]= 16'hd438;
assign i[7385]= 16'hd843;
assign i[7386]= 16'hdcf9;
assign i[7387]= 16'he247;
assign i[7388]= 16'he818;
assign i[7389]= 16'hee4e;
assign i[7390]= 16'hf4c9;
assign i[7391]= 16'hfb64;
assign i[7392]= 16'h1f8;
assign i[7393]= 16'h85f;
assign i[7394]= 16'he71;
assign i[7395]= 16'h1407;
assign i[7396]= 16'h1900;
assign i[7397]= 16'h1d3a;
assign i[7398]= 16'h209a;
assign i[7399]= 16'h230d;
assign i[7400]= 16'h2481;
assign i[7401]= 16'h24ef;
assign i[7402]= 16'h2453;
assign i[7403]= 16'h22b2;
assign i[7404]= 16'h2016;
assign i[7405]= 16'h1c90;
assign i[7406]= 16'h1836;
assign i[7407]= 16'h1321;
assign i[7408]= 16'hd70;
assign i[7409]= 16'h742;
assign i[7410]= 16'hbb;
assign i[7411]= 16'hf9fe;
assign i[7412]= 16'hf32d;
assign i[7413]= 16'hec6a;
assign i[7414]= 16'he5d7;
assign i[7415]= 16'hdf91;
assign i[7416]= 16'hd9b4;
assign i[7417]= 16'hd457;
assign i[7418]= 16'hcf8e;
assign i[7419]= 16'hcb6b;
assign i[7420]= 16'hc7f9;
assign i[7421]= 16'hc540;
assign i[7422]= 16'hc346;
assign i[7423]= 16'hc20d;
assign i[7424]= 16'hc190;
assign i[7425]= 16'hc1cd;
assign i[7426]= 16'hc2b9;
assign i[7427]= 16'hc44d;
assign i[7428]= 16'hc67a;
assign i[7429]= 16'hc933;
assign i[7430]= 16'hcc69;
assign i[7431]= 16'hd009;
assign i[7432]= 16'hd403;
assign i[7433]= 16'hd844;
assign i[7434]= 16'hdcb8;
assign i[7435]= 16'he14d;
assign i[7436]= 16'he5ee;
assign i[7437]= 16'hea89;
assign i[7438]= 16'hef0a;
assign i[7439]= 16'hf360;
assign i[7440]= 16'hf779;
assign i[7441]= 16'hfb44;
assign i[7442]= 16'hfeb4;
assign i[7443]= 16'h1bb;
assign i[7444]= 16'h450;
assign i[7445]= 16'h66a;
assign i[7446]= 16'h803;
assign i[7447]= 16'h918;
assign i[7448]= 16'h9ab;
assign i[7449]= 16'h9be;
assign i[7450]= 16'h958;
assign i[7451]= 16'h882;
assign i[7452]= 16'h74a;
assign i[7453]= 16'h5be;
assign i[7454]= 16'h3f1;
assign i[7455]= 16'h1f6;
assign i[7456]= 16'hffe3;
assign i[7457]= 16'hfdcc;
assign i[7458]= 16'hfbca;
assign i[7459]= 16'hf9f1;
assign i[7460]= 16'hf857;
assign i[7461]= 16'hf711;
assign i[7462]= 16'hf62e;
assign i[7463]= 16'hf5be;
assign i[7464]= 16'hf5cd;
assign i[7465]= 16'hf661;
assign i[7466]= 16'hf781;
assign i[7467]= 16'hf92a;
assign i[7468]= 16'hfb5a;
assign i[7469]= 16'hfe09;
assign i[7470]= 16'h128;
assign i[7471]= 16'h4ac;
assign i[7472]= 16'h881;
assign i[7473]= 16'hc92;
assign i[7474]= 16'h10c8;
assign i[7475]= 16'h150b;
assign i[7476]= 16'h1943;
assign i[7477]= 16'h1d56;
assign i[7478]= 16'h212e;
assign i[7479]= 16'h24b2;
assign i[7480]= 16'h27cf;
assign i[7481]= 16'h2a72;
assign i[7482]= 16'h2c8c;
assign i[7483]= 16'h2e11;
assign i[7484]= 16'h2ef8;
assign i[7485]= 16'h2f3c;
assign i[7486]= 16'h2edc;
assign i[7487]= 16'h2dda;
assign i[7488]= 16'h2c3a;
assign i[7489]= 16'h2a06;
assign i[7490]= 16'h2748;
assign i[7491]= 16'h240e;
assign i[7492]= 16'h2066;
assign i[7493]= 16'h1c62;
assign i[7494]= 16'h1814;
assign i[7495]= 16'h138c;
assign i[7496]= 16'hede;
assign i[7497]= 16'ha1b;
assign i[7498]= 16'h554;
assign i[7499]= 16'h9a;
assign i[7500]= 16'hfbfb;
assign i[7501]= 16'hf783;
assign i[7502]= 16'hf33f;
assign i[7503]= 16'hef39;
assign i[7504]= 16'heb79;
assign i[7505]= 16'he805;
assign i[7506]= 16'he4e2;
assign i[7507]= 16'he215;
assign i[7508]= 16'hdfa0;
assign i[7509]= 16'hdd83;
assign i[7510]= 16'hdbc0;
assign i[7511]= 16'hda54;
assign i[7512]= 16'hd941;
assign i[7513]= 16'hd883;
assign i[7514]= 16'hd819;
assign i[7515]= 16'hd800;
assign i[7516]= 16'hd835;
assign i[7517]= 16'hd8b7;
assign i[7518]= 16'hd980;
assign i[7519]= 16'hda8e;
assign i[7520]= 16'hdbdc;
assign i[7521]= 16'hdd66;
assign i[7522]= 16'hdf26;
assign i[7523]= 16'he117;
assign i[7524]= 16'he331;
assign i[7525]= 16'he56d;
assign i[7526]= 16'he7c1;
assign i[7527]= 16'hea25;
assign i[7528]= 16'hec8d;
assign i[7529]= 16'heeee;
assign i[7530]= 16'hf13c;
assign i[7531]= 16'hf369;
assign i[7532]= 16'hf56a;
assign i[7533]= 16'hf730;
assign i[7534]= 16'hf8b0;
assign i[7535]= 16'hf9de;
assign i[7536]= 16'hfaae;
assign i[7537]= 16'hfb17;
assign i[7538]= 16'hfb13;
assign i[7539]= 16'hfa9c;
assign i[7540]= 16'hf9b0;
assign i[7541]= 16'hf84f;
assign i[7542]= 16'hf67e;
assign i[7543]= 16'hf443;
assign i[7544]= 16'hf1aa;
assign i[7545]= 16'heebf;
assign i[7546]= 16'heb94;
assign i[7547]= 16'he83c;
assign i[7548]= 16'he4cf;
assign i[7549]= 16'he163;
assign i[7550]= 16'hde12;
assign i[7551]= 16'hdaf7;
assign i[7552]= 16'hd82c;
assign i[7553]= 16'hd5c9;
assign i[7554]= 16'hd3e7;
assign i[7555]= 16'hd29b;
assign i[7556]= 16'hd1f7;
assign i[7557]= 16'hd208;
assign i[7558]= 16'hd2da;
assign i[7559]= 16'hd471;
assign i[7560]= 16'hd6ce;
assign i[7561]= 16'hd9eb;
assign i[7562]= 16'hddbd;
assign i[7563]= 16'he235;
assign i[7564]= 16'he73f;
assign i[7565]= 16'hecc3;
assign i[7566]= 16'hf2a4;
assign i[7567]= 16'hf8c3;
assign i[7568]= 16'hff00;
assign i[7569]= 16'h538;
assign i[7570]= 16'hb4b;
assign i[7571]= 16'h1119;
assign i[7572]= 16'h1683;
assign i[7573]= 16'h1b6d;
assign i[7574]= 16'h1fc0;
assign i[7575]= 16'h236a;
assign i[7576]= 16'h265c;
assign i[7577]= 16'h288f;
assign i[7578]= 16'h2a00;
assign i[7579]= 16'h2ab2;
assign i[7580]= 16'h2aae;
assign i[7581]= 16'h2a02;
assign i[7582]= 16'h28c0;
assign i[7583]= 16'h2700;
assign i[7584]= 16'h24da;
assign i[7585]= 16'h226a;
assign i[7586]= 16'h1fcd;
assign i[7587]= 16'h1d20;
assign i[7588]= 16'h1a80;
assign i[7589]= 16'h1808;
assign i[7590]= 16'h15d0;
assign i[7591]= 16'h13ed;
assign i[7592]= 16'h1270;
assign i[7593]= 16'h1167;
assign i[7594]= 16'h10da;
assign i[7595]= 16'h10cc;
assign i[7596]= 16'h113d;
assign i[7597]= 16'h1227;
assign i[7598]= 16'h1382;
assign i[7599]= 16'h1540;
assign i[7600]= 16'h1751;
assign i[7601]= 16'h19a3;
assign i[7602]= 16'h1c22;
assign i[7603]= 16'h1eb8;
assign i[7604]= 16'h2151;
assign i[7605]= 16'h23d7;
assign i[7606]= 16'h2637;
assign i[7607]= 16'h285d;
assign i[7608]= 16'h2a3a;
assign i[7609]= 16'h2bbe;
assign i[7610]= 16'h2cde;
assign i[7611]= 16'h2d90;
assign i[7612]= 16'h2dce;
assign i[7613]= 16'h2d93;
assign i[7614]= 16'h2cde;
assign i[7615]= 16'h2bb0;
assign i[7616]= 16'h2a0a;
assign i[7617]= 16'h27f2;
assign i[7618]= 16'h256d;
assign i[7619]= 16'h2284;
assign i[7620]= 16'h1f3d;
assign i[7621]= 16'h1ba4;
assign i[7622]= 16'h17c1;
assign i[7623]= 16'h13a1;
assign i[7624]= 16'hf4e;
assign i[7625]= 16'had4;
assign i[7626]= 16'h63f;
assign i[7627]= 16'h19d;
assign i[7628]= 16'hfcfa;
assign i[7629]= 16'hf864;
assign i[7630]= 16'hf3e7;
assign i[7631]= 16'hef92;
assign i[7632]= 16'heb73;
assign i[7633]= 16'he796;
assign i[7634]= 16'he408;
assign i[7635]= 16'he0d6;
assign i[7636]= 16'hde0a;
assign i[7637]= 16'hdbad;
assign i[7638]= 16'hd9c8;
assign i[7639]= 16'hd85f;
assign i[7640]= 16'hd776;
assign i[7641]= 16'hd70c;
assign i[7642]= 16'hd721;
assign i[7643]= 16'hd7ad;
assign i[7644]= 16'hd8a8;
assign i[7645]= 16'hda06;
assign i[7646]= 16'hdbba;
assign i[7647]= 16'hddb2;
assign i[7648]= 16'hdfdb;
assign i[7649]= 16'he220;
assign i[7650]= 16'he46e;
assign i[7651]= 16'he6ad;
assign i[7652]= 16'he8c8;
assign i[7653]= 16'heaac;
assign i[7654]= 16'hec46;
assign i[7655]= 16'hed87;
assign i[7656]= 16'hee61;
assign i[7657]= 16'heecd;
assign i[7658]= 16'heec3;
assign i[7659]= 16'hee45;
assign i[7660]= 16'hed53;
assign i[7661]= 16'hebf6;
assign i[7662]= 16'hea39;
assign i[7663]= 16'he829;
assign i[7664]= 16'he5d8;
assign i[7665]= 16'he358;
assign i[7666]= 16'he0be;
assign i[7667]= 16'hde20;
assign i[7668]= 16'hdb90;
assign i[7669]= 16'hd924;
assign i[7670]= 16'hd6ec;
assign i[7671]= 16'hd4f7;
assign i[7672]= 16'hd351;
assign i[7673]= 16'hd201;
assign i[7674]= 16'hd10b;
assign i[7675]= 16'hd070;
assign i[7676]= 16'hd02a;
assign i[7677]= 16'hd032;
assign i[7678]= 16'hd07d;
assign i[7679]= 16'hd0fc;
assign i[7680]= 16'hd1a1;
assign i[7681]= 16'hd258;
assign i[7682]= 16'hd311;
assign i[7683]= 16'hd3bb;
assign i[7684]= 16'hd445;
assign i[7685]= 16'hd4a3;
assign i[7686]= 16'hd4c9;
assign i[7687]= 16'hd4b1;
assign i[7688]= 16'hd458;
assign i[7689]= 16'hd3be;
assign i[7690]= 16'hd2e8;
assign i[7691]= 16'hd1e2;
assign i[7692]= 16'hd0b8;
assign i[7693]= 16'hcf7b;
assign i[7694]= 16'hce3f;
assign i[7695]= 16'hcd1a;
assign i[7696]= 16'hcc24;
assign i[7697]= 16'hcb73;
assign i[7698]= 16'hcb1f;
assign i[7699]= 16'hcb3d;
assign i[7700]= 16'hcbe0;
assign i[7701]= 16'hcd16;
assign i[7702]= 16'hceeb;
assign i[7703]= 16'hd166;
assign i[7704]= 16'hd489;
assign i[7705]= 16'hd84f;
assign i[7706]= 16'hdcb0;
assign i[7707]= 16'he19e;
assign i[7708]= 16'he706;
assign i[7709]= 16'hecd2;
assign i[7710]= 16'hf2e7;
assign i[7711]= 16'hf928;
assign i[7712]= 16'hff75;
assign i[7713]= 16'h5ae;
assign i[7714]= 16'hbb4;
assign i[7715]= 16'h1167;
assign i[7716]= 16'h16a9;
assign i[7717]= 16'h1b60;
assign i[7718]= 16'h1f72;
assign i[7719]= 16'h22cd;
assign i[7720]= 16'h2560;
assign i[7721]= 16'h2722;
assign i[7722]= 16'h280b;
assign i[7723]= 16'h281a;
assign i[7724]= 16'h2754;
assign i[7725]= 16'h25c0;
assign i[7726]= 16'h236b;
assign i[7727]= 16'h2064;
assign i[7728]= 16'h1cbf;
assign i[7729]= 16'h1890;
assign i[7730]= 16'h13f0;
assign i[7731]= 16'hef8;
assign i[7732]= 16'h9c0;
assign i[7733]= 16'h463;
assign i[7734]= 16'hfef9;
assign i[7735]= 16'hf99a;
assign i[7736]= 16'hf45b;
assign i[7737]= 16'hef52;
assign i[7738]= 16'hea90;
assign i[7739]= 16'he627;
assign i[7740]= 16'he222;
assign i[7741]= 16'hde8e;
assign i[7742]= 16'hdb71;
assign i[7743]= 16'hd8d3;
assign i[7744]= 16'hd6b7;
assign i[7745]= 16'hd51e;
assign i[7746]= 16'hd407;
assign i[7747]= 16'hd370;
assign i[7748]= 16'hd355;
assign i[7749]= 16'hd3b0;
assign i[7750]= 16'hd47c;
assign i[7751]= 16'hd5b2;
assign i[7752]= 16'hd748;
assign i[7753]= 16'hd938;
assign i[7754]= 16'hdb78;
assign i[7755]= 16'hddff;
assign i[7756]= 16'he0c6;
assign i[7757]= 16'he3c4;
assign i[7758]= 16'he6ef;
assign i[7759]= 16'hea3f;
assign i[7760]= 16'hedad;
assign i[7761]= 16'hf12f;
assign i[7762]= 16'hf4be;
assign i[7763]= 16'hf853;
assign i[7764]= 16'hfbe4;
assign i[7765]= 16'hff69;
assign i[7766]= 16'h2da;
assign i[7767]= 16'h630;
assign i[7768]= 16'h962;
assign i[7769]= 16'hc66;
assign i[7770]= 16'hf34;
assign i[7771]= 16'h11c3;
assign i[7772]= 16'h1409;
assign i[7773]= 16'h15fd;
assign i[7774]= 16'h1797;
assign i[7775]= 16'h18ce;
assign i[7776]= 16'h199a;
assign i[7777]= 16'h19f4;
assign i[7778]= 16'h19d7;
assign i[7779]= 16'h193e;
assign i[7780]= 16'h1826;
assign i[7781]= 16'h1690;
assign i[7782]= 16'h147d;
assign i[7783]= 16'h11f1;
assign i[7784]= 16'hef3;
assign i[7785]= 16'hb8b;
assign i[7786]= 16'h7c7;
assign i[7787]= 16'h3b5;
assign i[7788]= 16'hff66;
assign i[7789]= 16'hfaeb;
assign i[7790]= 16'hf65b;
assign i[7791]= 16'hf1ca;
assign i[7792]= 16'hed51;
assign i[7793]= 16'he904;
assign i[7794]= 16'he4fb;
assign i[7795]= 16'he14a;
assign i[7796]= 16'hde05;
assign i[7797]= 16'hdb3b;
assign i[7798]= 16'hd8fb;
assign i[7799]= 16'hd74e;
assign i[7800]= 16'hd639;
assign i[7801]= 16'hd5be;
assign i[7802]= 16'hd5db;
assign i[7803]= 16'hd686;
assign i[7804]= 16'hd7b6;
assign i[7805]= 16'hd959;
assign i[7806]= 16'hdb5e;
assign i[7807]= 16'hddad;
assign i[7808]= 16'he030;
assign i[7809]= 16'he2cc;
assign i[7810]= 16'he56a;
assign i[7811]= 16'he7ef;
assign i[7812]= 16'hea46;
assign i[7813]= 16'hec5a;
assign i[7814]= 16'hee1b;
assign i[7815]= 16'hef7b;
assign i[7816]= 16'hf074;
assign i[7817]= 16'hf102;
assign i[7818]= 16'hf127;
assign i[7819]= 16'hf0ed;
assign i[7820]= 16'hf060;
assign i[7821]= 16'hef91;
assign i[7822]= 16'hee96;
assign i[7823]= 16'hed88;
assign i[7824]= 16'hec81;
assign i[7825]= 16'heb9d;
assign i[7826]= 16'heaf8;
assign i[7827]= 16'heaab;
assign i[7828]= 16'heacf;
assign i[7829]= 16'heb77;
assign i[7830]= 16'hecb2;
assign i[7831]= 16'hee8a;
assign i[7832]= 16'hf103;
assign i[7833]= 16'hf418;
assign i[7834]= 16'hf7c1;
assign i[7835]= 16'hfbed;
assign i[7836]= 16'h84;
assign i[7837]= 16'h56c;
assign i[7838]= 16'ha83;
assign i[7839]= 16'hfa5;
assign i[7840]= 16'h14a9;
assign i[7841]= 16'h1969;
assign i[7842]= 16'h1dbc;
assign i[7843]= 16'h217d;
assign i[7844]= 16'h2489;
assign i[7845]= 16'h26c2;
assign i[7846]= 16'h2810;
assign i[7847]= 16'h2862;
assign i[7848]= 16'h27ae;
assign i[7849]= 16'h25f2;
assign i[7850]= 16'h2336;
assign i[7851]= 16'h1f87;
assign i[7852]= 16'h1afe;
assign i[7853]= 16'h15b8;
assign i[7854]= 16'hfd9;
assign i[7855]= 16'h98b;
assign i[7856]= 16'h2fc;
assign i[7857]= 16'hfc5d;
assign i[7858]= 16'hf5de;
assign i[7859]= 16'hefaf;
assign i[7860]= 16'he9ff;
assign i[7861]= 16'he4fa;
assign i[7862]= 16'he0c6;
assign i[7863]= 16'hdd82;
assign i[7864]= 16'hdb48;
assign i[7865]= 16'hda29;
assign i[7866]= 16'hda2f;
assign i[7867]= 16'hdb5b;
assign i[7868]= 16'hdda7;
assign i[7869]= 16'he103;
assign i[7870]= 16'he55a;
assign i[7871]= 16'hea90;
assign i[7872]= 16'hf083;
assign i[7873]= 16'hf70d;
assign i[7874]= 16'hfe05;
assign i[7875]= 16'h541;
assign i[7876]= 16'hc98;
assign i[7877]= 16'h13de;
assign i[7878]= 16'h1aeb;
assign i[7879]= 16'h219a;
assign i[7880]= 16'h27cb;
assign i[7881]= 16'h2d61;
assign i[7882]= 16'h3244;
assign i[7883]= 16'h3663;
assign i[7884]= 16'h39b2;
assign i[7885]= 16'h3c2a;
assign i[7886]= 16'h3dc9;
assign i[7887]= 16'h3e93;
assign i[7888]= 16'h3e90;
assign i[7889]= 16'h3dcc;
assign i[7890]= 16'h3c54;
assign i[7891]= 16'h3a3a;
assign i[7892]= 16'h378f;
assign i[7893]= 16'h3466;
assign i[7894]= 16'h30d3;
assign i[7895]= 16'h2ce6;
assign i[7896]= 16'h28b0;
assign i[7897]= 16'h2441;
assign i[7898]= 16'h1fa7;
assign i[7899]= 16'h1aeb;
assign i[7900]= 16'h1618;
assign i[7901]= 16'h1135;
assign i[7902]= 16'hc47;
assign i[7903]= 16'h753;
assign i[7904]= 16'h25b;
assign i[7905]= 16'hfd63;
assign i[7906]= 16'hf86b;
assign i[7907]= 16'hf377;
assign i[7908]= 16'hee8a;
assign i[7909]= 16'he9a9;
assign i[7910]= 16'he4d9;
assign i[7911]= 16'he023;
assign i[7912]= 16'hdb91;
assign i[7913]= 16'hd72d;
assign i[7914]= 16'hd306;
assign i[7915]= 16'hcf2a;
assign i[7916]= 16'hcbaa;
assign i[7917]= 16'hc898;
assign i[7918]= 16'hc606;
assign i[7919]= 16'hc404;
assign i[7920]= 16'hc2a4;
assign i[7921]= 16'hc1f4;
assign i[7922]= 16'hc203;
assign i[7923]= 16'hc2d9;
assign i[7924]= 16'hc47e;
assign i[7925]= 16'hc6f3;
assign i[7926]= 16'hca37;
assign i[7927]= 16'hce43;
assign i[7928]= 16'hd309;
assign i[7929]= 16'hd87a;
assign i[7930]= 16'hde7f;
assign i[7931]= 16'he4fe;
assign i[7932]= 16'hebd6;
assign i[7933]= 16'hf2e7;
assign i[7934]= 16'hfa0a;
assign i[7935]= 16'h117;
assign i[7936]= 16'h7e9;
assign i[7937]= 16'he56;
assign i[7938]= 16'h1439;
assign i[7939]= 16'h196e;
assign i[7940]= 16'h1dd5;
assign i[7941]= 16'h2151;
assign i[7942]= 16'h23ce;
assign i[7943]= 16'h253b;
assign i[7944]= 16'h2590;
assign i[7945]= 16'h24cb;
assign i[7946]= 16'h22f2;
assign i[7947]= 16'h2012;
assign i[7948]= 16'h1c40;
assign i[7949]= 16'h1797;
assign i[7950]= 16'h1237;
assign i[7951]= 16'hc47;
assign i[7952]= 16'h5f0;
assign i[7953]= 16'hff5e;
assign i[7954]= 16'hf8bd;
assign i[7955]= 16'hf23a;
assign i[7956]= 16'hec00;
assign i[7957]= 16'he638;
assign i[7958]= 16'he104;
assign i[7959]= 16'hdc84;
assign i[7960]= 16'hd8ce;
assign i[7961]= 16'hd5f5;
assign i[7962]= 16'hd400;
assign i[7963]= 16'hd2f3;
assign i[7964]= 16'hd2c5;
assign i[7965]= 16'hd36b;
assign i[7966]= 16'hd4d0;
assign i[7967]= 16'hd6da;
assign i[7968]= 16'hd96c;
assign i[7969]= 16'hdc62;
assign i[7970]= 16'hdf99;
assign i[7971]= 16'he2ec;
assign i[7972]= 16'he638;
assign i[7973]= 16'he95c;
assign i[7974]= 16'hec38;
assign i[7975]= 16'heeb4;
assign i[7976]= 16'hf0bd;
assign i[7977]= 16'hf246;
assign i[7978]= 16'hf348;
assign i[7979]= 16'hf3c5;
assign i[7980]= 16'hf3c4;
assign i[7981]= 16'hf355;
assign i[7982]= 16'hf28b;
assign i[7983]= 16'hf181;
assign i[7984]= 16'hf053;
assign i[7985]= 16'hef20;
assign i[7986]= 16'hee0a;
assign i[7987]= 16'hed31;
assign i[7988]= 16'hecb3;
assign i[7989]= 16'hecab;
assign i[7990]= 16'hed2f;
assign i[7991]= 16'hee50;
assign i[7992]= 16'hf018;
assign i[7993]= 16'hf28b;
assign i[7994]= 16'hf5a3;
assign i[7995]= 16'hf954;
assign i[7996]= 16'hfd8d;
assign i[7997]= 16'h232;
assign i[7998]= 16'h727;
assign i[7999]= 16'hc47;
assign i[8000]= 16'h116c;
assign i[8001]= 16'h166d;
assign i[8002]= 16'h1b23;
assign i[8003]= 16'h1f66;
assign i[8004]= 16'h2314;
assign i[8005]= 16'h260d;
assign i[8006]= 16'h2838;
assign i[8007]= 16'h2982;
assign i[8008]= 16'h29e1;
assign i[8009]= 16'h2952;
assign i[8010]= 16'h27d9;
assign i[8011]= 16'h2586;
assign i[8012]= 16'h226d;
assign i[8013]= 16'h1eaa;
assign i[8014]= 16'h1a5f;
assign i[8015]= 16'h15b4;
assign i[8016]= 16'h10d3;
assign i[8017]= 16'hbe7;
assign i[8018]= 16'h71c;
assign i[8019]= 16'h29e;
assign i[8020]= 16'hfe95;
assign i[8021]= 16'hfb22;
assign i[8022]= 16'hf864;
assign i[8023]= 16'hf673;
assign i[8024]= 16'hf55d;
assign i[8025]= 16'hf52c;
assign i[8026]= 16'hf5e0;
assign i[8027]= 16'hf770;
assign i[8028]= 16'hf9ce;
assign i[8029]= 16'hfce4;
assign i[8030]= 16'h96;
assign i[8031]= 16'h4c4;
assign i[8032]= 16'h94b;
assign i[8033]= 16'he05;
assign i[8034]= 16'h12cc;
assign i[8035]= 16'h1778;
assign i[8036]= 16'h1be8;
assign i[8037]= 16'h1ffa;
assign i[8038]= 16'h2393;
assign i[8039]= 16'h269b;
assign i[8040]= 16'h2900;
assign i[8041]= 16'h2ab9;
assign i[8042]= 16'h2bbf;
assign i[8043]= 16'h2c15;
assign i[8044]= 16'h2bc1;
assign i[8045]= 16'h2ad1;
assign i[8046]= 16'h2956;
assign i[8047]= 16'h2765;
assign i[8048]= 16'h2518;
assign i[8049]= 16'h2288;
assign i[8050]= 16'h1fd2;
assign i[8051]= 16'h1d11;
assign i[8052]= 16'h1a60;
assign i[8053]= 16'h17d8;
assign i[8054]= 16'h158f;
assign i[8055]= 16'h1398;
assign i[8056]= 16'h1205;
assign i[8057]= 16'h10e0;
assign i[8058]= 16'h1031;
assign i[8059]= 16'hffd;
assign i[8060]= 16'h1044;
assign i[8061]= 16'h1103;
assign i[8062]= 16'h1231;
assign i[8063]= 16'h13c7;
assign i[8064]= 16'h15b9;
assign i[8065]= 16'h17f8;
assign i[8066]= 16'h1a76;
assign i[8067]= 16'h1d23;
assign i[8068]= 16'h1fef;
assign i[8069]= 16'h22ca;
assign i[8070]= 16'h25a5;
assign i[8071]= 16'h2870;
assign i[8072]= 16'h2b1e;
assign i[8073]= 16'h2da2;
assign i[8074]= 16'h2ff0;
assign i[8075]= 16'h31fd;
assign i[8076]= 16'h33c1;
assign i[8077]= 16'h3533;
assign i[8078]= 16'h364c;
assign i[8079]= 16'h3707;
assign i[8080]= 16'h375f;
assign i[8081]= 16'h3750;
assign i[8082]= 16'h36d8;
assign i[8083]= 16'h35f7;
assign i[8084]= 16'h34ac;
assign i[8085]= 16'h32f8;
assign i[8086]= 16'h30de;
assign i[8087]= 16'h2e63;
assign i[8088]= 16'h2b8d;
assign i[8089]= 16'h2863;
assign i[8090]= 16'h24ef;
assign i[8091]= 16'h213b;
assign i[8092]= 16'h1d54;
assign i[8093]= 16'h1949;
assign i[8094]= 16'h1528;
assign i[8095]= 16'h1104;
assign i[8096]= 16'hcec;
assign i[8097]= 16'h8f4;
assign i[8098]= 16'h52c;
assign i[8099]= 16'h1a6;
assign i[8100]= 16'hfe73;
assign i[8101]= 16'hfba0;
assign i[8102]= 16'hf93b;
assign i[8103]= 16'hf74f;
assign i[8104]= 16'hf5e3;
assign i[8105]= 16'hf4fb;
assign i[8106]= 16'hf498;
assign i[8107]= 16'hf4b9;
assign i[8108]= 16'hf556;
assign i[8109]= 16'hf667;
assign i[8110]= 16'hf7e0;
assign i[8111]= 16'hf9af;
assign i[8112]= 16'hfbc4;
assign i[8113]= 16'hfe0a;
assign i[8114]= 16'h6c;
assign i[8115]= 16'h2d4;
assign i[8116]= 16'h52c;
assign i[8117]= 16'h75f;
assign i[8118]= 16'h958;
assign i[8119]= 16'hb07;
assign i[8120]= 16'hc5a;
assign i[8121]= 16'hd46;
assign i[8122]= 16'hdc2;
assign i[8123]= 16'hdc9;
assign i[8124]= 16'hd58;
assign i[8125]= 16'hc71;
assign i[8126]= 16'hb1b;
assign i[8127]= 16'h95d;
assign i[8128]= 16'h743;
assign i[8129]= 16'h4db;
assign i[8130]= 16'h235;
assign i[8131]= 16'hff61;
assign i[8132]= 16'hfc6e;
assign i[8133]= 16'hf96f;
assign i[8134]= 16'hf673;
assign i[8135]= 16'hf389;
assign i[8136]= 16'hf0bb;
assign i[8137]= 16'hee16;
assign i[8138]= 16'heb9e;
assign i[8139]= 16'he95a;
assign i[8140]= 16'he74b;
assign i[8141]= 16'he56f;
assign i[8142]= 16'he3c2;
assign i[8143]= 16'he240;
assign i[8144]= 16'he0df;
assign i[8145]= 16'hdf97;
assign i[8146]= 16'hde5f;
assign i[8147]= 16'hdd2e;
assign i[8148]= 16'hdbfa;
assign i[8149]= 16'hdabb;
assign i[8150]= 16'hd96d;
assign i[8151]= 16'hd80b;
assign i[8152]= 16'hd694;
assign i[8153]= 16'hd50a;
assign i[8154]= 16'hd372;
assign i[8155]= 16'hd1d4;
assign i[8156]= 16'hd039;
assign i[8157]= 16'hceae;
assign i[8158]= 16'hcd43;
assign i[8159]= 16'hcc07;
assign i[8160]= 16'hcb0a;
assign i[8161]= 16'hca5e;
assign i[8162]= 16'hca12;
assign i[8163]= 16'hca36;
assign i[8164]= 16'hcad5;
assign i[8165]= 16'hcbf8;
assign i[8166]= 16'hcda6;
assign i[8167]= 16'hcfe1;
assign i[8168]= 16'hd2a5;
assign i[8169]= 16'hd5eb;
assign i[8170]= 16'hd9a8;
assign i[8171]= 16'hddcc;
assign i[8172]= 16'he242;
assign i[8173]= 16'he6f2;
assign i[8174]= 16'hebc3;
assign i[8175]= 16'hf096;
assign i[8176]= 16'hf54e;
assign i[8177]= 16'hf9cc;
assign i[8178]= 16'hfdf3;
assign i[8179]= 16'h1a4;
assign i[8180]= 16'h4c9;
assign i[8181]= 16'h74b;
assign i[8182]= 16'h918;
assign i[8183]= 16'ha23;
assign i[8184]= 16'ha65;
assign i[8185]= 16'h9dd;
assign i[8186]= 16'h890;
assign i[8187]= 16'h688;
assign i[8188]= 16'h3d5;
assign i[8189]= 16'h8c;
assign i[8190]= 16'hfcc8;
assign i[8191]= 16'hf8a3;
assign i[8192]= 16'hf43f;
assign i[8193]= 16'hefbd;
assign i[8194]= 16'heb3d;
assign i[8195]= 16'he6e2;
assign i[8196]= 16'he2cb;
assign i[8197]= 16'hdf14;
assign i[8198]= 16'hdbd5;
assign i[8199]= 16'hd924;
assign i[8200]= 16'hd710;
assign i[8201]= 16'hd5a2;
assign i[8202]= 16'hd4df;
assign i[8203]= 16'hd4c4;
assign i[8204]= 16'hd549;
assign i[8205]= 16'hd663;
assign i[8206]= 16'hd7ff;
assign i[8207]= 16'hda08;
assign i[8208]= 16'hdc65;
assign i[8209]= 16'hdefc;
assign i[8210]= 16'he1b0;
assign i[8211]= 16'he466;
assign i[8212]= 16'he701;
assign i[8213]= 16'he968;
assign i[8214]= 16'heb85;
assign i[8215]= 16'hed44;
assign i[8216]= 16'hee94;
assign i[8217]= 16'hef6b;
assign i[8218]= 16'hefc2;
assign i[8219]= 16'hef97;
assign i[8220]= 16'heeed;
assign i[8221]= 16'hedca;
assign i[8222]= 16'hec3a;
assign i[8223]= 16'hea4b;
assign i[8224]= 16'he80c;
assign i[8225]= 16'he591;
assign i[8226]= 16'he2ed;
assign i[8227]= 16'he035;
assign i[8228]= 16'hdd7c;
assign i[8229]= 16'hdad4;
assign i[8230]= 16'hd84e;
assign i[8231]= 16'hd5fa;
assign i[8232]= 16'hd3e2;
assign i[8233]= 16'hd211;
assign i[8234]= 16'hd08c;
assign i[8235]= 16'hcf56;
assign i[8236]= 16'hce70;
assign i[8237]= 16'hcdd8;
assign i[8238]= 16'hcd8a;
assign i[8239]= 16'hcd7f;
assign i[8240]= 16'hcdb1;
assign i[8241]= 16'hce17;
assign i[8242]= 16'hcea9;
assign i[8243]= 16'hcf5f;
assign i[8244]= 16'hd030;
assign i[8245]= 16'hd118;
assign i[8246]= 16'hd20f;
assign i[8247]= 16'hd313;
assign i[8248]= 16'hd420;
assign i[8249]= 16'hd537;
assign i[8250]= 16'hd657;
assign i[8251]= 16'hd783;
assign i[8252]= 16'hd8bd;
assign i[8253]= 16'hda09;
assign i[8254]= 16'hdb6c;
assign i[8255]= 16'hdcea;
assign i[8256]= 16'hde87;
assign i[8257]= 16'he049;
assign i[8258]= 16'he231;
assign i[8259]= 16'he443;
assign i[8260]= 16'he680;
assign i[8261]= 16'he8e9;
assign i[8262]= 16'heb7e;
assign i[8263]= 16'hee3d;
assign i[8264]= 16'hf124;
assign i[8265]= 16'hf430;
assign i[8266]= 16'hf75d;
assign i[8267]= 16'hfaa7;
assign i[8268]= 16'hfe0a;
assign i[8269]= 16'h181;
assign i[8270]= 16'h508;
assign i[8271]= 16'h89b;
assign i[8272]= 16'hc35;
assign i[8273]= 16'hfd3;
assign i[8274]= 16'h1370;
assign i[8275]= 16'h1709;
assign i[8276]= 16'h1a99;
assign i[8277]= 16'h1e1b;
assign i[8278]= 16'h218c;
assign i[8279]= 16'h24e5;
assign i[8280]= 16'h2820;
assign i[8281]= 16'h2b36;
assign i[8282]= 16'h2e1c;
assign i[8283]= 16'h30cb;
assign i[8284]= 16'h3338;
assign i[8285]= 16'h3556;
assign i[8286]= 16'h371a;
assign i[8287]= 16'h3876;
assign i[8288]= 16'h395f;
assign i[8289]= 16'h39c8;
assign i[8290]= 16'h39a7;
assign i[8291]= 16'h38f1;
assign i[8292]= 16'h379f;
assign i[8293]= 16'h35ac;
assign i[8294]= 16'h3316;
assign i[8295]= 16'h2fde;
assign i[8296]= 16'h2c09;
assign i[8297]= 16'h27a0;
assign i[8298]= 16'h22b0;
assign i[8299]= 16'h1d48;
assign i[8300]= 16'h177e;
assign i[8301]= 16'h1167;
assign i[8302]= 16'hb1d;
assign i[8303]= 16'h4bd;
assign i[8304]= 16'hfe63;
assign i[8305]= 16'hf82c;
assign i[8306]= 16'hf234;
assign i[8307]= 16'hec97;
assign i[8308]= 16'he76f;
assign i[8309]= 16'he2d1;
assign i[8310]= 16'hded0;
assign i[8311]= 16'hdb7b;
assign i[8312]= 16'hd8db;
assign i[8313]= 16'hd6f5;
assign i[8314]= 16'hd5c8;
assign i[8315]= 16'hd550;
assign i[8316]= 16'hd581;
assign i[8317]= 16'hd64f;
assign i[8318]= 16'hd7a6;
assign i[8319]= 16'hd971;
assign i[8320]= 16'hdb9a;
assign i[8321]= 16'hde08;
assign i[8322]= 16'he0a2;
assign i[8323]= 16'he34e;
assign i[8324]= 16'he5f6;
assign i[8325]= 16'he885;
assign i[8326]= 16'heae7;
assign i[8327]= 16'hed0d;
assign i[8328]= 16'heeec;
assign i[8329]= 16'hf07b;
assign i[8330]= 16'hf1b7;
assign i[8331]= 16'hf2a0;
assign i[8332]= 16'hf339;
assign i[8333]= 16'hf38a;
assign i[8334]= 16'hf39c;
assign i[8335]= 16'hf37b;
assign i[8336]= 16'hf335;
assign i[8337]= 16'hf2d8;
assign i[8338]= 16'hf273;
assign i[8339]= 16'hf214;
assign i[8340]= 16'hf1c9;
assign i[8341]= 16'hf19e;
assign i[8342]= 16'hf19e;
assign i[8343]= 16'hf1cf;
assign i[8344]= 16'hf239;
assign i[8345]= 16'hf2dd;
assign i[8346]= 16'hf3bd;
assign i[8347]= 16'hf4d8;
assign i[8348]= 16'hf628;
assign i[8349]= 16'hf7aa;
assign i[8350]= 16'hf955;
assign i[8351]= 16'hfb22;
assign i[8352]= 16'hfd06;
assign i[8353]= 16'hfef8;
assign i[8354]= 16'hee;
assign i[8355]= 16'h2de;
assign i[8356]= 16'h4bd;
assign i[8357]= 16'h683;
assign i[8358]= 16'h826;
assign i[8359]= 16'h99e;
assign i[8360]= 16'hae2;
assign i[8361]= 16'hbea;
assign i[8362]= 16'hcb1;
assign i[8363]= 16'hd30;
assign i[8364]= 16'hd61;
assign i[8365]= 16'hd3e;
assign i[8366]= 16'hcc3;
assign i[8367]= 16'hbec;
assign i[8368]= 16'hab6;
assign i[8369]= 16'h91f;
assign i[8370]= 16'h725;
assign i[8371]= 16'h4c9;
assign i[8372]= 16'h20e;
assign i[8373]= 16'hfefa;
assign i[8374]= 16'hfb90;
assign i[8375]= 16'hf7dc;
assign i[8376]= 16'hf3ea;
assign i[8377]= 16'hefc8;
assign i[8378]= 16'heb89;
assign i[8379]= 16'he740;
assign i[8380]= 16'he303;
assign i[8381]= 16'hdeec;
assign i[8382]= 16'hdb13;
assign i[8383]= 16'hd793;
assign i[8384]= 16'hd487;
assign i[8385]= 16'hd208;
assign i[8386]= 16'hd02e;
assign i[8387]= 16'hcf0d;
assign i[8388]= 16'hceb7;
assign i[8389]= 16'hcf3a;
assign i[8390]= 16'hd09c;
assign i[8391]= 16'hd2e0;
assign i[8392]= 16'hd603;
assign i[8393]= 16'hd9f9;
assign i[8394]= 16'hdeb2;
assign i[8395]= 16'he417;
assign i[8396]= 16'hea0b;
assign i[8397]= 16'hf06c;
assign i[8398]= 16'hf712;
assign i[8399]= 16'hfdd5;
assign i[8400]= 16'h488;
assign i[8401]= 16'haff;
assign i[8402]= 16'h110f;
assign i[8403]= 16'h168c;
assign i[8404]= 16'h1b50;
assign i[8405]= 16'h1f39;
assign i[8406]= 16'h222b;
assign i[8407]= 16'h2410;
assign i[8408]= 16'h24db;
assign i[8409]= 16'h2486;
assign i[8410]= 16'h2314;
assign i[8411]= 16'h208f;
assign i[8412]= 16'h1d0a;
assign i[8413]= 16'h18a1;
assign i[8414]= 16'h1374;
assign i[8415]= 16'hda9;
assign i[8416]= 16'h76c;
assign i[8417]= 16'heb;
assign i[8418]= 16'hfa56;
assign i[8419]= 16'hf3db;
assign i[8420]= 16'heda9;
assign i[8421]= 16'he7ec;
assign i[8422]= 16'he2ca;
assign i[8423]= 16'hde65;
assign i[8424]= 16'hdada;
assign i[8425]= 16'hd83d;
assign i[8426]= 16'hd69d;
assign i[8427]= 16'hd600;
assign i[8428]= 16'hd664;
assign i[8429]= 16'hd7c3;
assign i[8430]= 16'hda0d;
assign i[8431]= 16'hdd2f;
assign i[8432]= 16'he10e;
assign i[8433]= 16'he58f;
assign i[8434]= 16'hea92;
assign i[8435]= 16'heff5;
assign i[8436]= 16'hf596;
assign i[8437]= 16'hfb55;
assign i[8438]= 16'h110;
assign i[8439]= 16'h6ac;
assign i[8440]= 16'hc0d;
assign i[8441]= 16'h111f;
assign i[8442]= 16'h15cd;
assign i[8443]= 16'h1a0b;
assign i[8444]= 16'h1dce;
assign i[8445]= 16'h2112;
assign i[8446]= 16'h23d6;
assign i[8447]= 16'h261c;
assign i[8448]= 16'h27e9;
assign i[8449]= 16'h2948;
assign i[8450]= 16'h2a43;
assign i[8451]= 16'h2ae5;
assign i[8452]= 16'h2b3d;
assign i[8453]= 16'h2b59;
assign i[8454]= 16'h2b45;
assign i[8455]= 16'h2b11;
assign i[8456]= 16'h2ac6;
assign i[8457]= 16'h2a73;
assign i[8458]= 16'h2a1f;
assign i[8459]= 16'h29d4;
assign i[8460]= 16'h2998;
assign i[8461]= 16'h2971;
assign i[8462]= 16'h2963;
assign i[8463]= 16'h2970;
assign i[8464]= 16'h299a;
assign i[8465]= 16'h29e1;
assign i[8466]= 16'h2a44;
assign i[8467]= 16'h2ac1;
assign i[8468]= 16'h2b57;
assign i[8469]= 16'h2c02;
assign i[8470]= 16'h2cbe;
assign i[8471]= 16'h2d87;
assign i[8472]= 16'h2e58;
assign i[8473]= 16'h2f2d;
assign i[8474]= 16'h2fff;
assign i[8475]= 16'h30c7;
assign i[8476]= 16'h317f;
assign i[8477]= 16'h321f;
assign i[8478]= 16'h329f;
assign i[8479]= 16'h32f7;
assign i[8480]= 16'h331e;
assign i[8481]= 16'h330b;
assign i[8482]= 16'h32b4;
assign i[8483]= 16'h3212;
assign i[8484]= 16'h311c;
assign i[8485]= 16'h2fca;
assign i[8486]= 16'h2e16;
assign i[8487]= 16'h2bfa;
assign i[8488]= 16'h2972;
assign i[8489]= 16'h267d;
assign i[8490]= 16'h2319;
assign i[8491]= 16'h1f4a;
assign i[8492]= 16'h1b12;
assign i[8493]= 16'h1678;
assign i[8494]= 16'h1185;
assign i[8495]= 16'hc44;
assign i[8496]= 16'h6c1;
assign i[8497]= 16'h10c;
assign i[8498]= 16'hfb35;
assign i[8499]= 16'hf54d;
assign i[8500]= 16'hef68;
assign i[8501]= 16'he998;
assign i[8502]= 16'he3f2;
assign i[8503]= 16'hde89;
assign i[8504]= 16'hd970;
assign i[8505]= 16'hd4b8;
assign i[8506]= 16'hd074;
assign i[8507]= 16'hccb2;
assign i[8508]= 16'hc97f;
assign i[8509]= 16'hc6e7;
assign i[8510]= 16'hc4f3;
assign i[8511]= 16'hc3a9;
assign i[8512]= 16'hc30d;
assign i[8513]= 16'hc321;
assign i[8514]= 16'hc3e5;
assign i[8515]= 16'hc554;
assign i[8516]= 16'hc769;
assign i[8517]= 16'hca1d;
assign i[8518]= 16'hcd64;
assign i[8519]= 16'hd135;
assign i[8520]= 16'hd580;
assign i[8521]= 16'hda37;
assign i[8522]= 16'hdf4b;
assign i[8523]= 16'he4a9;
assign i[8524]= 16'hea40;
assign i[8525]= 16'heffe;
assign i[8526]= 16'hf5cf;
assign i[8527]= 16'hfba2;
assign i[8528]= 16'h162;
assign i[8529]= 16'h700;
assign i[8530]= 16'hc68;
assign i[8531]= 16'h118b;
assign i[8532]= 16'h1658;
assign i[8533]= 16'h1ac2;
assign i[8534]= 16'h1ebb;
assign i[8535]= 16'h2239;
assign i[8536]= 16'h2533;
assign i[8537]= 16'h27a1;
assign i[8538]= 16'h297e;
assign i[8539]= 16'h2ac8;
assign i[8540]= 16'h2b7e;
assign i[8541]= 16'h2ba2;
assign i[8542]= 16'h2b38;
assign i[8543]= 16'h2a45;
assign i[8544]= 16'h28d3;
assign i[8545]= 16'h26eb;
assign i[8546]= 16'h249a;
assign i[8547]= 16'h21ec;
assign i[8548]= 16'h1ef0;
assign i[8549]= 16'h1bb6;
assign i[8550]= 16'h184d;
assign i[8551]= 16'h14c7;
assign i[8552]= 16'h1132;
assign i[8553]= 16'hda0;
assign i[8554]= 16'ha1f;
assign i[8555]= 16'h6be;
assign i[8556]= 16'h389;
assign i[8557]= 16'h8b;
assign i[8558]= 16'hfdd1;
assign i[8559]= 16'hfb5f;
assign i[8560]= 16'hf93e;
assign i[8561]= 16'hf771;
assign i[8562]= 16'hf5fc;
assign i[8563]= 16'hf4df;
assign i[8564]= 16'hf419;
assign i[8565]= 16'hf3a8;
assign i[8566]= 16'hf389;
assign i[8567]= 16'hf3b7;
assign i[8568]= 16'hf42b;
assign i[8569]= 16'hf4e1;
assign i[8570]= 16'hf5d0;
assign i[8571]= 16'hf6f2;
assign i[8572]= 16'hf83e;
assign i[8573]= 16'hf9af;
assign i[8574]= 16'hfb3d;
assign i[8575]= 16'hfce0;
assign i[8576]= 16'hfe93;
assign i[8577]= 16'h4f;
assign i[8578]= 16'h20f;
assign i[8579]= 16'h3ce;
assign i[8580]= 16'h587;
assign i[8581]= 16'h736;
assign i[8582]= 16'h8d6;
assign i[8583]= 16'ha64;
assign i[8584]= 16'hbdc;
assign i[8585]= 16'hd3b;
assign i[8586]= 16'he7d;
assign i[8587]= 16'hfa1;
assign i[8588]= 16'h10a3;
assign i[8589]= 16'h117f;
assign i[8590]= 16'h1235;
assign i[8591]= 16'h12c2;
assign i[8592]= 16'h1325;
assign i[8593]= 16'h135b;
assign i[8594]= 16'h1366;
assign i[8595]= 16'h1345;
assign i[8596]= 16'h12f9;
assign i[8597]= 16'h1285;
assign i[8598]= 16'h11ec;
assign i[8599]= 16'h1132;
assign i[8600]= 16'h105c;
assign i[8601]= 16'hf72;
assign i[8602]= 16'he7a;
assign i[8603]= 16'hd7e;
assign i[8604]= 16'hc87;
assign i[8605]= 16'hb9e;
assign i[8606]= 16'hace;
assign i[8607]= 16'ha20;
assign i[8608]= 16'h9a0;
assign i[8609]= 16'h956;
assign i[8610]= 16'h94b;
assign i[8611]= 16'h985;
assign i[8612]= 16'ha0b;
assign i[8613]= 16'hae0;
assign i[8614]= 16'hc04;
assign i[8615]= 16'hd78;
assign i[8616]= 16'hf38;
assign i[8617]= 16'h113d;
assign i[8618]= 16'h137e;
assign i[8619]= 16'h15f1;
assign i[8620]= 16'h1888;
assign i[8621]= 16'h1b32;
assign i[8622]= 16'h1de0;
assign i[8623]= 16'h207e;
assign i[8624]= 16'h22f9;
assign i[8625]= 16'h253f;
assign i[8626]= 16'h273c;
assign i[8627]= 16'h28df;
assign i[8628]= 16'h2a18;
assign i[8629]= 16'h2ad8;
assign i[8630]= 16'h2b15;
assign i[8631]= 16'h2ac7;
assign i[8632]= 16'h29e9;
assign i[8633]= 16'h287b;
assign i[8634]= 16'h2680;
assign i[8635]= 16'h23ff;
assign i[8636]= 16'h2104;
assign i[8637]= 16'h1d9f;
assign i[8638]= 16'h19e0;
assign i[8639]= 16'h15dc;
assign i[8640]= 16'h11ac;
assign i[8641]= 16'hd67;
assign i[8642]= 16'h928;
assign i[8643]= 16'h507;
assign i[8644]= 16'h11d;
assign i[8645]= 16'hfd83;
assign i[8646]= 16'hfa4c;
assign i[8647]= 16'hf78b;
assign i[8648]= 16'hf54f;
assign i[8649]= 16'hf3a3;
assign i[8650]= 16'hf28e;
assign i[8651]= 16'hf213;
assign i[8652]= 16'hf22f;
assign i[8653]= 16'hf2de;
assign i[8654]= 16'hf416;
assign i[8655]= 16'hf5ca;
assign i[8656]= 16'hf7ea;
assign i[8657]= 16'hfa64;
assign i[8658]= 16'hfd25;
assign i[8659]= 16'h18;
assign i[8660]= 16'h329;
assign i[8661]= 16'h646;
assign i[8662]= 16'h95c;
assign i[8663]= 16'hc5a;
assign i[8664]= 16'hf35;
assign i[8665]= 16'h11e1;
assign i[8666]= 16'h1457;
assign i[8667]= 16'h1695;
assign i[8668]= 16'h1899;
assign i[8669]= 16'h1a67;
assign i[8670]= 16'h1c03;
assign i[8671]= 16'h1d76;
assign i[8672]= 16'h1ec9;
assign i[8673]= 16'h2007;
assign i[8674]= 16'h213c;
assign i[8675]= 16'h2270;
assign i[8676]= 16'h23b0;
assign i[8677]= 16'h2501;
assign i[8678]= 16'h266b;
assign i[8679]= 16'h27f0;
assign i[8680]= 16'h298f;
assign i[8681]= 16'h2b47;
assign i[8682]= 16'h2d0f;
assign i[8683]= 16'h2ede;
assign i[8684]= 16'h30a7;
assign i[8685]= 16'h325a;
assign i[8686]= 16'h33e6;
assign i[8687]= 16'h3538;
assign i[8688]= 16'h363c;
assign i[8689]= 16'h36df;
assign i[8690]= 16'h370e;
assign i[8691]= 16'h36b9;
assign i[8692]= 16'h35d1;
assign i[8693]= 16'h344d;
assign i[8694]= 16'h3224;
assign i[8695]= 16'h2f54;
assign i[8696]= 16'h2bdf;
assign i[8697]= 16'h27cb;
assign i[8698]= 16'h2324;
assign i[8699]= 16'h1dfa;
assign i[8700]= 16'h1860;
assign i[8701]= 16'h126d;
assign i[8702]= 16'hc3d;
assign i[8703]= 16'h5eb;
assign i[8704]= 16'hff97;
assign i[8705]= 16'hf95d;
assign i[8706]= 16'hf35c;
assign i[8707]= 16'hedaf;
assign i[8708]= 16'he872;
assign i[8709]= 16'he3bb;
assign i[8710]= 16'hdf9e;
assign i[8711]= 16'hdc29;
assign i[8712]= 16'hd967;
assign i[8713]= 16'hd75e;
assign i[8714]= 16'hd60e;
assign i[8715]= 16'hd572;
assign i[8716]= 16'hd582;
assign i[8717]= 16'hd62f;
assign i[8718]= 16'hd768;
assign i[8719]= 16'hd919;
assign i[8720]= 16'hdb29;
assign i[8721]= 16'hdd81;
assign i[8722]= 16'he006;
assign i[8723]= 16'he29e;
assign i[8724]= 16'he52e;
assign i[8725]= 16'he7a0;
assign i[8726]= 16'he9dc;
assign i[8727]= 16'hebcf;
assign i[8728]= 16'hed67;
assign i[8729]= 16'hee98;
assign i[8730]= 16'hef57;
assign i[8731]= 16'hef9f;
assign i[8732]= 16'hef6d;
assign i[8733]= 16'heec3;
assign i[8734]= 16'heda6;
assign i[8735]= 16'hec1d;
assign i[8736]= 16'hea34;
assign i[8737]= 16'he7f7;
assign i[8738]= 16'he577;
assign i[8739]= 16'he2c3;
assign i[8740]= 16'hdfed;
assign i[8741]= 16'hdd07;
assign i[8742]= 16'hda22;
assign i[8743]= 16'hd74f;
assign i[8744]= 16'hd49f;
assign i[8745]= 16'hd220;
assign i[8746]= 16'hcfe0;
assign i[8747]= 16'hcdeb;
assign i[8748]= 16'hcc49;
assign i[8749]= 16'hcb02;
assign i[8750]= 16'hca1c;
assign i[8751]= 16'hc99a;
assign i[8752]= 16'hc97e;
assign i[8753]= 16'hc9c6;
assign i[8754]= 16'hca71;
assign i[8755]= 16'hcb7c;
assign i[8756]= 16'hcce1;
assign i[8757]= 16'hce9b;
assign i[8758]= 16'hd0a4;
assign i[8759]= 16'hd2f3;
assign i[8760]= 16'hd582;
assign i[8761]= 16'hd848;
assign i[8762]= 16'hdb3e;
assign i[8763]= 16'hde5d;
assign i[8764]= 16'he19d;
assign i[8765]= 16'he4f7;
assign i[8766]= 16'he863;
assign i[8767]= 16'hebdc;
assign i[8768]= 16'hef5b;
assign i[8769]= 16'hf2da;
assign i[8770]= 16'hf654;
assign i[8771]= 16'hf9c2;
assign i[8772]= 16'hfd1f;
assign i[8773]= 16'h64;
assign i[8774]= 16'h38e;
assign i[8775]= 16'h695;
assign i[8776]= 16'h973;
assign i[8777]= 16'hc22;
assign i[8778]= 16'he9a;
assign i[8779]= 16'h10d7;
assign i[8780]= 16'h12d0;
assign i[8781]= 16'h147f;
assign i[8782]= 16'h15df;
assign i[8783]= 16'h16e9;
assign i[8784]= 16'h179a;
assign i[8785]= 16'h17ed;
assign i[8786]= 16'h17df;
assign i[8787]= 16'h1770;
assign i[8788]= 16'h16a0;
assign i[8789]= 16'h1572;
assign i[8790]= 16'h13ea;
assign i[8791]= 16'h120e;
assign i[8792]= 16'hfe8;
assign i[8793]= 16'hd82;
assign i[8794]= 16'hae8;
assign i[8795]= 16'h828;
assign i[8796]= 16'h553;
assign i[8797]= 16'h279;
assign i[8798]= 16'hffab;
assign i[8799]= 16'hfcfa;
assign i[8800]= 16'hfa77;
assign i[8801]= 16'hf833;
assign i[8802]= 16'hf63c;
assign i[8803]= 16'hf4a0;
assign i[8804]= 16'hf369;
assign i[8805]= 16'hf29f;
assign i[8806]= 16'hf247;
assign i[8807]= 16'hf262;
assign i[8808]= 16'hf2ef;
assign i[8809]= 16'hf3e7;
assign i[8810]= 16'hf543;
assign i[8811]= 16'hf6f6;
assign i[8812]= 16'hf8f1;
assign i[8813]= 16'hfb23;
assign i[8814]= 16'hfd7a;
assign i[8815]= 16'hffe0;
assign i[8816]= 16'h241;
assign i[8817]= 16'h489;
assign i[8818]= 16'h6a3;
assign i[8819]= 16'h87e;
assign i[8820]= 16'ha09;
assign i[8821]= 16'hb36;
assign i[8822]= 16'hbfc;
assign i[8823]= 16'hc54;
assign i[8824]= 16'hc3b;
assign i[8825]= 16'hbb3;
assign i[8826]= 16'hac1;
assign i[8827]= 16'h96e;
assign i[8828]= 16'h7c7;
assign i[8829]= 16'h5db;
assign i[8830]= 16'h3bd;
assign i[8831]= 16'h182;
assign i[8832]= 16'hff3f;
assign i[8833]= 16'hfd08;
assign i[8834]= 16'hfaf6;
assign i[8835]= 16'hf91c;
assign i[8836]= 16'hf78f;
assign i[8837]= 16'hf660;
assign i[8838]= 16'hf59e;
assign i[8839]= 16'hf554;
assign i[8840]= 16'hf58c;
assign i[8841]= 16'hf648;
assign i[8842]= 16'hf78b;
assign i[8843]= 16'hf951;
assign i[8844]= 16'hfb95;
assign i[8845]= 16'hfe4c;
assign i[8846]= 16'h169;
assign i[8847]= 16'h4de;
assign i[8848]= 16'h89a;
assign i[8849]= 16'hc8a;
assign i[8850]= 16'h1098;
assign i[8851]= 16'h14b1;
assign i[8852]= 16'h18bf;
assign i[8853]= 16'h1caf;
assign i[8854]= 16'h206b;
assign i[8855]= 16'h23e1;
assign i[8856]= 16'h2701;
assign i[8857]= 16'h29b8;
assign i[8858]= 16'h2bfb;
assign i[8859]= 16'h2dbb;
assign i[8860]= 16'h2ef0;
assign i[8861]= 16'h2f92;
assign i[8862]= 16'h2f9a;
assign i[8863]= 16'h2f06;
assign i[8864]= 16'h2dd4;
assign i[8865]= 16'h2c05;
assign i[8866]= 16'h299c;
assign i[8867]= 16'h26a1;
assign i[8868]= 16'h2319;
assign i[8869]= 16'h1f11;
assign i[8870]= 16'h1a95;
assign i[8871]= 16'h15b3;
assign i[8872]= 16'h107e;
assign i[8873]= 16'hb08;
assign i[8874]= 16'h567;
assign i[8875]= 16'hffb2;
assign i[8876]= 16'hfa00;
assign i[8877]= 16'hf46c;
assign i[8878]= 16'hef0f;
assign i[8879]= 16'hea04;
assign i[8880]= 16'he564;
assign i[8881]= 16'he148;
assign i[8882]= 16'hddc7;
assign i[8883]= 16'hdaf5;
assign i[8884]= 16'hd8e5;
assign i[8885]= 16'hd7a4;
assign i[8886]= 16'hd73c;
assign i[8887]= 16'hd7b4;
assign i[8888]= 16'hd90b;
assign i[8889]= 16'hdb3d;
assign i[8890]= 16'hde40;
assign i[8891]= 16'he207;
assign i[8892]= 16'he67c;
assign i[8893]= 16'heb88;
assign i[8894]= 16'hf10f;
assign i[8895]= 16'hf6f2;
assign i[8896]= 16'hfd0e;
assign i[8897]= 16'h341;
assign i[8898]= 16'h968;
assign i[8899]= 16'hf5f;
assign i[8900]= 16'h1505;
assign i[8901]= 16'h1a3c;
assign i[8902]= 16'h1ee7;
assign i[8903]= 16'h22f1;
assign i[8904]= 16'h2648;
assign i[8905]= 16'h28de;
assign i[8906]= 16'h2aae;
assign i[8907]= 16'h2bb7;
assign i[8908]= 16'h2bff;
assign i[8909]= 16'h2b8f;
assign i[8910]= 16'h2a78;
assign i[8911]= 16'h28cf;
assign i[8912]= 16'h26aa;
assign i[8913]= 16'h2426;
assign i[8914]= 16'h215d;
assign i[8915]= 16'h1e6c;
assign i[8916]= 16'h1b71;
assign i[8917]= 16'h1885;
assign i[8918]= 16'h15c0;
assign i[8919]= 16'h1339;
assign i[8920]= 16'h1101;
assign i[8921]= 16'hf23;
assign i[8922]= 16'hda8;
assign i[8923]= 16'hc93;
assign i[8924]= 16'hbe2;
assign i[8925]= 16'hb8f;
assign i[8926]= 16'hb8e;
assign i[8927]= 16'hbd1;
assign i[8928]= 16'hc47;
assign i[8929]= 16'hcdc;
assign i[8930]= 16'hd7b;
assign i[8931]= 16'he0f;
assign i[8932]= 16'he81;
assign i[8933]= 16'hebf;
assign i[8934]= 16'heb6;
assign i[8935]= 16'he57;
assign i[8936]= 16'hd94;
assign i[8937]= 16'hc65;
assign i[8938]= 16'hac5;
assign i[8939]= 16'h8b2;
assign i[8940]= 16'h62d;
assign i[8941]= 16'h33d;
assign i[8942]= 16'hffec;
assign i[8943]= 16'hfc42;
assign i[8944]= 16'hf84f;
assign i[8945]= 16'hf423;
assign i[8946]= 16'hefcf;
assign i[8947]= 16'heb64;
assign i[8948]= 16'he6f6;
assign i[8949]= 16'he296;
assign i[8950]= 16'hde55;
assign i[8951]= 16'hda44;
assign i[8952]= 16'hd672;
assign i[8953]= 16'hd2ed;
assign i[8954]= 16'hcfc1;
assign i[8955]= 16'hccf9;
assign i[8956]= 16'hca9e;
assign i[8957]= 16'hc8b7;
assign i[8958]= 16'hc74c;
assign i[8959]= 16'hc661;
assign i[8960]= 16'hc5f8;
assign i[8961]= 16'hc616;
assign i[8962]= 16'hc6bb;
assign i[8963]= 16'hc7e8;
assign i[8964]= 16'hc99b;
assign i[8965]= 16'hcbd4;
assign i[8966]= 16'hce8e;
assign i[8967]= 16'hd1c6;
assign i[8968]= 16'hd576;
assign i[8969]= 16'hd997;
assign i[8970]= 16'hde1f;
assign i[8971]= 16'he305;
assign i[8972]= 16'he83c;
assign i[8973]= 16'hedb7;
assign i[8974]= 16'hf364;
assign i[8975]= 16'hf935;
assign i[8976]= 16'hff15;
assign i[8977]= 16'h4f2;
assign i[8978]= 16'haba;
assign i[8979]= 16'h1058;
assign i[8980]= 16'h15b9;
assign i[8981]= 16'h1aca;
assign i[8982]= 16'h1f7b;
assign i[8983]= 16'h23bd;
assign i[8984]= 16'h2784;
assign i[8985]= 16'h2ac8;
assign i[8986]= 16'h2d82;
assign i[8987]= 16'h2faf;
assign i[8988]= 16'h3153;
assign i[8989]= 16'h3271;
assign i[8990]= 16'h3312;
assign i[8991]= 16'h3342;
assign i[8992]= 16'h3311;
assign i[8993]= 16'h328f;
assign i[8994]= 16'h31cf;
assign i[8995]= 16'h30e4;
assign i[8996]= 16'h2fe2;
assign i[8997]= 16'h2edd;
assign i[8998]= 16'h2de6;
assign i[8999]= 16'h2d0d;
assign i[9000]= 16'h2c5f;
assign i[9001]= 16'h2be4;
assign i[9002]= 16'h2ba4;
assign i[9003]= 16'h2ba1;
assign i[9004]= 16'h2bd7;
assign i[9005]= 16'h2c41;
assign i[9006]= 16'h2cd6;
assign i[9007]= 16'h2d8a;
assign i[9008]= 16'h2e4c;
assign i[9009]= 16'h2f0c;
assign i[9010]= 16'h2fb8;
assign i[9011]= 16'h303e;
assign i[9012]= 16'h308c;
assign i[9013]= 16'h3094;
assign i[9014]= 16'h3048;
assign i[9015]= 16'h2f9f;
assign i[9016]= 16'h2e92;
assign i[9017]= 16'h2d21;
assign i[9018]= 16'h2b4e;
assign i[9019]= 16'h2922;
assign i[9020]= 16'h26a8;
assign i[9021]= 16'h23f1;
assign i[9022]= 16'h2110;
assign i[9023]= 16'h1e1e;
assign i[9024]= 16'h1b33;
assign i[9025]= 16'h1867;
assign i[9026]= 16'h15d7;
assign i[9027]= 16'h1399;
assign i[9028]= 16'h11c4;
assign i[9029]= 16'h106b;
assign i[9030]= 16'hf9d;
assign i[9031]= 16'hf63;
assign i[9032]= 16'hfc2;
assign i[9033]= 16'h10b8;
assign i[9034]= 16'h123d;
assign i[9035]= 16'h1442;
assign i[9036]= 16'h16b5;
assign i[9037]= 16'h197d;
assign i[9038]= 16'h1c7c;
assign i[9039]= 16'h1f92;
assign i[9040]= 16'h229d;
assign i[9041]= 16'h2578;
assign i[9042]= 16'h2801;
assign i[9043]= 16'h2a16;
assign i[9044]= 16'h2b98;
assign i[9045]= 16'h2c6c;
assign i[9046]= 16'h2c7d;
assign i[9047]= 16'h2bbb;
assign i[9048]= 16'h2a1e;
assign i[9049]= 16'h27a3;
assign i[9050]= 16'h2450;
assign i[9051]= 16'h2031;
assign i[9052]= 16'h1b59;
assign i[9053]= 16'h15e3;
assign i[9054]= 16'hfeb;
assign i[9055]= 16'h997;
assign i[9056]= 16'h30a;
assign i[9057]= 16'hfc6f;
assign i[9058]= 16'hf5eb;
assign i[9059]= 16'hefa7;
assign i[9060]= 16'he9c7;
assign i[9061]= 16'he46d;
assign i[9062]= 16'hdfb7;
assign i[9063]= 16'hdbba;
assign i[9064]= 16'hd888;
assign i[9065]= 16'hd62c;
assign i[9066]= 16'hd4a8;
assign i[9067]= 16'hd3fa;
assign i[9068]= 16'hd416;
assign i[9069]= 16'hd4ed;
assign i[9070]= 16'hd669;
assign i[9071]= 16'hd86e;
assign i[9072]= 16'hdae0;
assign i[9073]= 16'hdd9d;
assign i[9074]= 16'he085;
assign i[9075]= 16'he376;
assign i[9076]= 16'he650;
assign i[9077]= 16'he8f4;
assign i[9078]= 16'heb48;
assign i[9079]= 16'hed37;
assign i[9080]= 16'heead;
assign i[9081]= 16'hef9e;
assign i[9082]= 16'hf004;
assign i[9083]= 16'hefdc;
assign i[9084]= 16'hef2b;
assign i[9085]= 16'hedf8;
assign i[9086]= 16'hec51;
assign i[9087]= 16'hea46;
assign i[9088]= 16'he7eb;
assign i[9089]= 16'he554;
assign i[9090]= 16'he299;
assign i[9091]= 16'hdfd0;
assign i[9092]= 16'hdd0e;
assign i[9093]= 16'hda67;
assign i[9094]= 16'hd7ef;
assign i[9095]= 16'hd5b4;
assign i[9096]= 16'hd3c2;
assign i[9097]= 16'hd221;
assign i[9098]= 16'hd0d6;
assign i[9099]= 16'hcfe2;
assign i[9100]= 16'hcf42;
assign i[9101]= 16'hcef1;
assign i[9102]= 16'hcee6;
assign i[9103]= 16'hcf17;
assign i[9104]= 16'hcf77;
assign i[9105]= 16'hcff9;
assign i[9106]= 16'hd091;
assign i[9107]= 16'hd130;
assign i[9108]= 16'hd1ca;
assign i[9109]= 16'hd256;
assign i[9110]= 16'hd2c9;
assign i[9111]= 16'hd31c;
assign i[9112]= 16'hd34d;
assign i[9113]= 16'hd359;
assign i[9114]= 16'hd340;
assign i[9115]= 16'hd307;
assign i[9116]= 16'hd2b3;
assign i[9117]= 16'hd24c;
assign i[9118]= 16'hd1db;
assign i[9119]= 16'hd16a;
assign i[9120]= 16'hd104;
assign i[9121]= 16'hd0b7;
assign i[9122]= 16'hd08c;
assign i[9123]= 16'hd08f;
assign i[9124]= 16'hd0ca;
assign i[9125]= 16'hd147;
assign i[9126]= 16'hd20c;
assign i[9127]= 16'hd320;
assign i[9128]= 16'hd486;
assign i[9129]= 16'hd640;
assign i[9130]= 16'hd850;
assign i[9131]= 16'hdab2;
assign i[9132]= 16'hdd64;
assign i[9133]= 16'he062;
assign i[9134]= 16'he3a4;
assign i[9135]= 16'he725;
assign i[9136]= 16'headb;
assign i[9137]= 16'heebd;
assign i[9138]= 16'hf2c3;
assign i[9139]= 16'hf6e3;
assign i[9140]= 16'hfb13;
assign i[9141]= 16'hff48;
assign i[9142]= 16'h379;
assign i[9143]= 16'h79e;
assign i[9144]= 16'hbac;
assign i[9145]= 16'hf9c;
assign i[9146]= 16'h1363;
assign i[9147]= 16'h16fb;
assign i[9148]= 16'h1a5b;
assign i[9149]= 16'h1d7e;
assign i[9150]= 16'h205b;
assign i[9151]= 16'h22ed;
assign i[9152]= 16'h2530;
assign i[9153]= 16'h271e;
assign i[9154]= 16'h28b5;
assign i[9155]= 16'h29f2;
assign i[9156]= 16'h2ad3;
assign i[9157]= 16'h2b58;
assign i[9158]= 16'h2b82;
assign i[9159]= 16'h2b54;
assign i[9160]= 16'h2ad2;
assign i[9161]= 16'h2a00;
assign i[9162]= 16'h28e5;
assign i[9163]= 16'h278a;
assign i[9164]= 16'h25f7;
assign i[9165]= 16'h2436;
assign i[9166]= 16'h2252;
assign i[9167]= 16'h2057;
assign i[9168]= 16'h1e50;
assign i[9169]= 16'h1c49;
assign i[9170]= 16'h1a4e;
assign i[9171]= 16'h1869;
assign i[9172]= 16'h16a3;
assign i[9173]= 16'h1506;
assign i[9174]= 16'h1399;
assign i[9175]= 16'h125f;
assign i[9176]= 16'h115d;
assign i[9177]= 16'h1094;
assign i[9178]= 16'h1001;
assign i[9179]= 16'hfa2;
assign i[9180]= 16'hf72;
assign i[9181]= 16'hf69;
assign i[9182]= 16'hf7e;
assign i[9183]= 16'hfa6;
assign i[9184]= 16'hfd6;
assign i[9185]= 16'h1002;
assign i[9186]= 16'h101c;
assign i[9187]= 16'h1019;
assign i[9188]= 16'hfea;
assign i[9189]= 16'hf86;
assign i[9190]= 16'hee2;
assign i[9191]= 16'hdf4;
assign i[9192]= 16'hcb7;
assign i[9193]= 16'hb23;
assign i[9194]= 16'h938;
assign i[9195]= 16'h6f3;
assign i[9196]= 16'h457;
assign i[9197]= 16'h167;
assign i[9198]= 16'hfe2b;
assign i[9199]= 16'hfaa9;
assign i[9200]= 16'hf6eb;
assign i[9201]= 16'hf2fe;
assign i[9202]= 16'heeee;
assign i[9203]= 16'heac9;
assign i[9204]= 16'he69e;
assign i[9205]= 16'he27c;
assign i[9206]= 16'hde72;
assign i[9207]= 16'hda90;
assign i[9208]= 16'hd6e3;
assign i[9209]= 16'hd37b;
assign i[9210]= 16'hd064;
assign i[9211]= 16'hcda9;
assign i[9212]= 16'hcb56;
assign i[9213]= 16'hc973;
assign i[9214]= 16'hc809;
assign i[9215]= 16'hc71d;
assign i[9216]= 16'hc6b4;
assign i[9217]= 16'hc6d1;
assign i[9218]= 16'hc775;
assign i[9219]= 16'hc89f;
assign i[9220]= 16'hca4e;
assign i[9221]= 16'hcc7e;
assign i[9222]= 16'hcf2a;
assign i[9223]= 16'hd24d;
assign i[9224]= 16'hd5df;
assign i[9225]= 16'hd9d7;
assign i[9226]= 16'hde2d;
assign i[9227]= 16'he2d4;
assign i[9228]= 16'he7c3;
assign i[9229]= 16'heced;
assign i[9230]= 16'hf245;
assign i[9231]= 16'hf7bf;
assign i[9232]= 16'hfd4d;
assign i[9233]= 16'h2e0;
assign i[9234]= 16'h86d;
assign i[9235]= 16'hde4;
assign i[9236]= 16'h1339;
assign i[9237]= 16'h185f;
assign i[9238]= 16'h1d49;
assign i[9239]= 16'h21ea;
assign i[9240]= 16'h2638;
assign i[9241]= 16'h2a28;
assign i[9242]= 16'h2db1;
assign i[9243]= 16'h30cb;
assign i[9244]= 16'h336d;
assign i[9245]= 16'h3594;
assign i[9246]= 16'h373a;
assign i[9247]= 16'h385b;
assign i[9248]= 16'h38f8;
assign i[9249]= 16'h3910;
assign i[9250]= 16'h38a4;
assign i[9251]= 16'h37b7;
assign i[9252]= 16'h364f;
assign i[9253]= 16'h3471;
assign i[9254]= 16'h3226;
assign i[9255]= 16'h2f76;
assign i[9256]= 16'h2c6b;
assign i[9257]= 16'h2911;
assign i[9258]= 16'h2575;
assign i[9259]= 16'h21a3;
assign i[9260]= 16'h1da9;
assign i[9261]= 16'h1996;
assign i[9262]= 16'h1579;
assign i[9263]= 16'h115f;
assign i[9264]= 16'hd56;
assign i[9265]= 16'h96c;
assign i[9266]= 16'h5ae;
assign i[9267]= 16'h226;
assign i[9268]= 16'hfee0;
assign i[9269]= 16'hfbe3;
assign i[9270]= 16'hf935;
assign i[9271]= 16'hf6dc;
assign i[9272]= 16'hf4da;
assign i[9273]= 16'hf330;
assign i[9274]= 16'hf1db;
assign i[9275]= 16'hf0d8;
assign i[9276]= 16'hf021;
assign i[9277]= 16'hefae;
assign i[9278]= 16'hef76;
assign i[9279]= 16'hef6e;
assign i[9280]= 16'hef8a;
assign i[9281]= 16'hefbe;
assign i[9282]= 16'heffd;
assign i[9283]= 16'hf03a;
assign i[9284]= 16'hf069;
assign i[9285]= 16'hf07e;
assign i[9286]= 16'hf070;
assign i[9287]= 16'hf035;
assign i[9288]= 16'hefc7;
assign i[9289]= 16'hef20;
assign i[9290]= 16'hee3e;
assign i[9291]= 16'hed20;
assign i[9292]= 16'hebc7;
assign i[9293]= 16'hea38;
assign i[9294]= 16'he877;
assign i[9295]= 16'he68d;
assign i[9296]= 16'he482;
assign i[9297]= 16'he25f;
assign i[9298]= 16'he02f;
assign i[9299]= 16'hddfe;
assign i[9300]= 16'hdbd6;
assign i[9301]= 16'hd9c1;
assign i[9302]= 16'hd7c9;
assign i[9303]= 16'hd5f7;
assign i[9304]= 16'hd453;
assign i[9305]= 16'hd2e1;
assign i[9306]= 16'hd1a7;
assign i[9307]= 16'hd0a6;
assign i[9308]= 16'hcfe0;
assign i[9309]= 16'hcf54;
assign i[9310]= 16'hceff;
assign i[9311]= 16'hcee0;
assign i[9312]= 16'hcef0;
assign i[9313]= 16'hcf2c;
assign i[9314]= 16'hcf8e;
assign i[9315]= 16'hd011;
assign i[9316]= 16'hd0b0;
assign i[9317]= 16'hd167;
assign i[9318]= 16'hd231;
assign i[9319]= 16'hd30c;
assign i[9320]= 16'hd3f7;
assign i[9321]= 16'hd4f0;
assign i[9322]= 16'hd5f8;
assign i[9323]= 16'hd710;
assign i[9324]= 16'hd83b;
assign i[9325]= 16'hd97c;
assign i[9326]= 16'hdad7;
assign i[9327]= 16'hdc4f;
assign i[9328]= 16'hddea;
assign i[9329]= 16'hdfaa;
assign i[9330]= 16'he194;
assign i[9331]= 16'he3aa;
assign i[9332]= 16'he5ef;
assign i[9333]= 16'he863;
assign i[9334]= 16'heb08;
assign i[9335]= 16'heddd;
assign i[9336]= 16'hf0de;
assign i[9337]= 16'hf40a;
assign i[9338]= 16'hf75d;
assign i[9339]= 16'hfad1;
assign i[9340]= 16'hfe61;
assign i[9341]= 16'h206;
assign i[9342]= 16'h5bc;
assign i[9343]= 16'h97b;
assign i[9344]= 16'hd3d;
assign i[9345]= 16'h10fa;
assign i[9346]= 16'h14ac;
assign i[9347]= 16'h184c;
assign i[9348]= 16'h1bd5;
assign i[9349]= 16'h1f3f;
assign i[9350]= 16'h2287;
assign i[9351]= 16'h25a4;
assign i[9352]= 16'h2893;
assign i[9353]= 16'h2b4d;
assign i[9354]= 16'h2dcc;
assign i[9355]= 16'h300b;
assign i[9356]= 16'h3203;
assign i[9357]= 16'h33af;
assign i[9358]= 16'h3509;
assign i[9359]= 16'h360a;
assign i[9360]= 16'h36ac;
assign i[9361]= 16'h36eb;
assign i[9362]= 16'h36c2;
assign i[9363]= 16'h362d;
assign i[9364]= 16'h3529;
assign i[9365]= 16'h33b5;
assign i[9366]= 16'h31d2;
assign i[9367]= 16'h2f83;
assign i[9368]= 16'h2ccc;
assign i[9369]= 16'h29b5;
assign i[9370]= 16'h2645;
assign i[9371]= 16'h228a;
assign i[9372]= 16'h1e90;
assign i[9373]= 16'h1a67;
assign i[9374]= 16'h161f;
assign i[9375]= 16'h11cc;
assign i[9376]= 16'hd7f;
assign i[9377]= 16'h94b;
assign i[9378]= 16'h543;
assign i[9379]= 16'h178;
assign i[9380]= 16'hfdfb;
assign i[9381]= 16'hfad6;
assign i[9382]= 16'hf816;
assign i[9383]= 16'hf5c2;
assign i[9384]= 16'hf3dd;
assign i[9385]= 16'hf268;
assign i[9386]= 16'hf15f;
assign i[9387]= 16'hf0bc;
assign i[9388]= 16'hf072;
assign i[9389]= 16'hf076;
assign i[9390]= 16'hf0b6;
assign i[9391]= 16'hf120;
assign i[9392]= 16'hf1a0;
assign i[9393]= 16'hf223;
assign i[9394]= 16'hf295;
assign i[9395]= 16'hf2e3;
assign i[9396]= 16'hf2fc;
assign i[9397]= 16'hf2d2;
assign i[9398]= 16'hf25a;
assign i[9399]= 16'hf18c;
assign i[9400]= 16'hf065;
assign i[9401]= 16'heee6;
assign i[9402]= 16'hed14;
assign i[9403]= 16'heaf9;
assign i[9404]= 16'he8a2;
assign i[9405]= 16'he61f;
assign i[9406]= 16'he385;
assign i[9407]= 16'he0e9;
assign i[9408]= 16'hde64;
assign i[9409]= 16'hdc0c;
assign i[9410]= 16'hd9fa;
assign i[9411]= 16'hd845;
assign i[9412]= 16'hd702;
assign i[9413]= 16'hd644;
assign i[9414]= 16'hd61b;
assign i[9415]= 16'hd692;
assign i[9416]= 16'hd7b1;
assign i[9417]= 16'hd97d;
assign i[9418]= 16'hdbf6;
assign i[9419]= 16'hdf16;
assign i[9420]= 16'he2d5;
assign i[9421]= 16'he727;
assign i[9422]= 16'hebfc;
assign i[9423]= 16'hf142;
assign i[9424]= 16'hf6e6;
assign i[9425]= 16'hfccf;
assign i[9426]= 16'h2e7;
assign i[9427]= 16'h918;
assign i[9428]= 16'hf49;
assign i[9429]= 16'h1562;
assign i[9430]= 16'h1b4e;
assign i[9431]= 16'h20f8;
assign i[9432]= 16'h264b;
assign i[9433]= 16'h2b37;
assign i[9434]= 16'h2fab;
assign i[9435]= 16'h3399;
assign i[9436]= 16'h36f6;
assign i[9437]= 16'h39b6;
assign i[9438]= 16'h3bd3;
assign i[9439]= 16'h3d44;
assign i[9440]= 16'h3e07;
assign i[9441]= 16'h3e17;
assign i[9442]= 16'h3d75;
assign i[9443]= 16'h3c20;
assign i[9444]= 16'h3a1d;
assign i[9445]= 16'h376f;
assign i[9446]= 16'h341e;
assign i[9447]= 16'h3034;
assign i[9448]= 16'h2bbb;
assign i[9449]= 16'h26c2;
assign i[9450]= 16'h2158;
assign i[9451]= 16'h1b91;
assign i[9452]= 16'h1580;
assign i[9453]= 16'hf3d;
assign i[9454]= 16'h8df;
assign i[9455]= 16'h280;
assign i[9456]= 16'hfc3b;
assign i[9457]= 16'hf628;
assign i[9458]= 16'hf061;
assign i[9459]= 16'heb00;
assign i[9460]= 16'he61a;
assign i[9461]= 16'he1c5;
assign i[9462]= 16'hde10;
assign i[9463]= 16'hdb09;
assign i[9464]= 16'hd8b8;
assign i[9465]= 16'hd721;
assign i[9466]= 16'hd643;
assign i[9467]= 16'hd619;
assign i[9468]= 16'hd696;
assign i[9469]= 16'hd7ad;
assign i[9470]= 16'hd949;
assign i[9471]= 16'hdb53;
assign i[9472]= 16'hddb1;
assign i[9473]= 16'he048;
assign i[9474]= 16'he2fc;
assign i[9475]= 16'he5b0;
assign i[9476]= 16'he84a;
assign i[9477]= 16'heab2;
assign i[9478]= 16'hecd2;
assign i[9479]= 16'hee9a;
assign i[9480]= 16'heffe;
assign i[9481]= 16'hf0f8;
assign i[9482]= 16'hf185;
assign i[9483]= 16'hf1ab;
assign i[9484]= 16'hf174;
assign i[9485]= 16'hf0f0;
assign i[9486]= 16'hf030;
assign i[9487]= 16'hef4d;
assign i[9488]= 16'hee61;
assign i[9489]= 16'hed86;
assign i[9490]= 16'hecd7;
assign i[9491]= 16'hec70;
assign i[9492]= 16'hec68;
assign i[9493]= 16'hecd4;
assign i[9494]= 16'hedc5;
assign i[9495]= 16'hef47;
assign i[9496]= 16'hf15f;
assign i[9497]= 16'hf40d;
assign i[9498]= 16'hf74a;
assign i[9499]= 16'hfb09;
assign i[9500]= 16'hff36;
assign i[9501]= 16'h3b8;
assign i[9502]= 16'h875;
assign i[9503]= 16'hd4a;
assign i[9504]= 16'h1214;
assign i[9505]= 16'h16af;
assign i[9506]= 16'h1af7;
assign i[9507]= 16'h1ec9;
assign i[9508]= 16'h2204;
assign i[9509]= 16'h248c;
assign i[9510]= 16'h2649;
assign i[9511]= 16'h2729;
assign i[9512]= 16'h271f;
assign i[9513]= 16'h2627;
assign i[9514]= 16'h2442;
assign i[9515]= 16'h2176;
assign i[9516]= 16'h1dd4;
assign i[9517]= 16'h196f;
assign i[9518]= 16'h1461;
assign i[9519]= 16'hec7;
assign i[9520]= 16'h8c2;
assign i[9521]= 16'h275;
assign i[9522]= 16'hfc07;
assign i[9523]= 16'hf599;
assign i[9524]= 16'hef50;
assign i[9525]= 16'he94f;
assign i[9526]= 16'he3b3;
assign i[9527]= 16'hde9a;
assign i[9528]= 16'hda1a;
assign i[9529]= 16'hd647;
assign i[9530]= 16'hd330;
assign i[9531]= 16'hd0de;
assign i[9532]= 16'hcf57;
assign i[9533]= 16'hce9d;
assign i[9534]= 16'hceac;
assign i[9535]= 16'hcf7e;
assign i[9536]= 16'hd109;
assign i[9537]= 16'hd340;
assign i[9538]= 16'hd614;
assign i[9539]= 16'hd976;
assign i[9540]= 16'hdd53;
assign i[9541]= 16'he199;
assign i[9542]= 16'he634;
assign i[9543]= 16'heb13;
assign i[9544]= 16'hf021;
assign i[9545]= 16'hf54d;
assign i[9546]= 16'hfa83;
assign i[9547]= 16'hffb4;
assign i[9548]= 16'h4cc;
assign i[9549]= 16'h9be;
assign i[9550]= 16'he7a;
assign i[9551]= 16'h12f1;
assign i[9552]= 16'h1717;
assign i[9553]= 16'h1adf;
assign i[9554]= 16'h1e40;
assign i[9555]= 16'h212f;
assign i[9556]= 16'h23a7;
assign i[9557]= 16'h25a1;
assign i[9558]= 16'h2719;
assign i[9559]= 16'h2811;
assign i[9560]= 16'h2888;
assign i[9561]= 16'h2883;
assign i[9562]= 16'h2809;
assign i[9563]= 16'h2723;
assign i[9564]= 16'h25dd;
assign i[9565]= 16'h2446;
assign i[9566]= 16'h226e;
assign i[9567]= 16'h2067;
assign i[9568]= 16'h1e44;
assign i[9569]= 16'h1c19;
assign i[9570]= 16'h19fb;
assign i[9571]= 16'h17fd;
assign i[9572]= 16'h1632;
assign i[9573]= 16'h14ab;
assign i[9574]= 16'h1376;
assign i[9575]= 16'h129f;
assign i[9576]= 16'h122e;
assign i[9577]= 16'h1228;
assign i[9578]= 16'h128f;
assign i[9579]= 16'h135f;
assign i[9580]= 16'h1491;
assign i[9581]= 16'h161d;
assign i[9582]= 16'h17f3;
assign i[9583]= 16'h1a04;
assign i[9584]= 16'h1c3d;
assign i[9585]= 16'h1e8b;
assign i[9586]= 16'h20d9;
assign i[9587]= 16'h2311;
assign i[9588]= 16'h251f;
assign i[9589]= 16'h26f2;
assign i[9590]= 16'h2878;
assign i[9591]= 16'h29a4;
assign i[9592]= 16'h2a6b;
assign i[9593]= 16'h2ac5;
assign i[9594]= 16'h2ab1;
assign i[9595]= 16'h2a2f;
assign i[9596]= 16'h2942;
assign i[9597]= 16'h27f4;
assign i[9598]= 16'h264f;
assign i[9599]= 16'h2463;
assign i[9600]= 16'h223f;
assign i[9601]= 16'h1ff6;
assign i[9602]= 16'h1d9c;
assign i[9603]= 16'h1b44;
assign i[9604]= 16'h1901;
assign i[9605]= 16'h16e7;
assign i[9606]= 16'h1505;
assign i[9607]= 16'h136c;
assign i[9608]= 16'h1228;
assign i[9609]= 16'h1142;
assign i[9610]= 16'h10c2;
assign i[9611]= 16'h10ac;
assign i[9612]= 16'h1101;
assign i[9613]= 16'h11c0;
assign i[9614]= 16'h12e3;
assign i[9615]= 16'h1465;
assign i[9616]= 16'h163b;
assign i[9617]= 16'h185d;
assign i[9618]= 16'h1abc;
assign i[9619]= 16'h1d4e;
assign i[9620]= 16'h2002;
assign i[9621]= 16'h22cc;
assign i[9622]= 16'h259e;
assign i[9623]= 16'h2868;
assign i[9624]= 16'h2b1d;
assign i[9625]= 16'h2db0;
assign i[9626]= 16'h3015;
assign i[9627]= 16'h323e;
assign i[9628]= 16'h3422;
assign i[9629]= 16'h35b5;
assign i[9630]= 16'h36ef;
assign i[9631]= 16'h37c6;
assign i[9632]= 16'h3832;
assign i[9633]= 16'h382d;
assign i[9634]= 16'h37b2;
assign i[9635]= 16'h36bc;
assign i[9636]= 16'h3547;
assign i[9637]= 16'h3352;
assign i[9638]= 16'h30de;
assign i[9639]= 16'h2deb;
assign i[9640]= 16'h2a7d;
assign i[9641]= 16'h269a;
assign i[9642]= 16'h224a;
assign i[9643]= 16'h1d95;
assign i[9644]= 16'h1889;
assign i[9645]= 16'h1331;
assign i[9646]= 16'hd9e;
assign i[9647]= 16'h7e0;
assign i[9648]= 16'h20a;
assign i[9649]= 16'hfc30;
assign i[9650]= 16'hf662;
assign i[9651]= 16'hf0b6;
assign i[9652]= 16'heb3d;
assign i[9653]= 16'he60b;
assign i[9654]= 16'he12f;
assign i[9655]= 16'hdcb8;
assign i[9656]= 16'hd8b2;
assign i[9657]= 16'hd527;
assign i[9658]= 16'hd21e;
assign i[9659]= 16'hcf9a;
assign i[9660]= 16'hcd9e;
assign i[9661]= 16'hcc25;
assign i[9662]= 16'hcb2d;
assign i[9663]= 16'hcaad;
assign i[9664]= 16'hca9c;
assign i[9665]= 16'hcaee;
assign i[9666]= 16'hcb98;
assign i[9667]= 16'hcc8b;
assign i[9668]= 16'hcdba;
assign i[9669]= 16'hcf19;
assign i[9670]= 16'hd099;
assign i[9671]= 16'hd231;
assign i[9672]= 16'hd3d5;
assign i[9673]= 16'hd57f;
assign i[9674]= 16'hd727;
assign i[9675]= 16'hd8ca;
assign i[9676]= 16'hda66;
assign i[9677]= 16'hdbfa;
assign i[9678]= 16'hdd88;
assign i[9679]= 16'hdf13;
assign i[9680]= 16'he09f;
assign i[9681]= 16'he231;
assign i[9682]= 16'he3cd;
assign i[9683]= 16'he57a;
assign i[9684]= 16'he73b;
assign i[9685]= 16'he913;
assign i[9686]= 16'heb06;
assign i[9687]= 16'hed13;
assign i[9688]= 16'hef3b;
assign i[9689]= 16'hf17b;
assign i[9690]= 16'hf3cf;
assign i[9691]= 16'hf632;
assign i[9692]= 16'hf89d;
assign i[9693]= 16'hfb08;
assign i[9694]= 16'hfd6b;
assign i[9695]= 16'hffbc;
assign i[9696]= 16'h1f1;
assign i[9697]= 16'h402;
assign i[9698]= 16'h5e5;
assign i[9699]= 16'h793;
assign i[9700]= 16'h905;
assign i[9701]= 16'ha34;
assign i[9702]= 16'hb1c;
assign i[9703]= 16'hbbb;
assign i[9704]= 16'hc0e;
assign i[9705]= 16'hc16;
assign i[9706]= 16'hbd4;
assign i[9707]= 16'hb4a;
assign i[9708]= 16'ha7b;
assign i[9709]= 16'h96d;
assign i[9710]= 16'h825;
assign i[9711]= 16'h6a7;
assign i[9712]= 16'h4fa;
assign i[9713]= 16'h325;
assign i[9714]= 16'h12e;
assign i[9715]= 16'hff1c;
assign i[9716]= 16'hfcf4;
assign i[9717]= 16'hfabe;
assign i[9718]= 16'hf882;
assign i[9719]= 16'hf646;
assign i[9720]= 16'hf412;
assign i[9721]= 16'hf1ee;
assign i[9722]= 16'hefe3;
assign i[9723]= 16'hedfa;
assign i[9724]= 16'hec3c;
assign i[9725]= 16'heab3;
assign i[9726]= 16'he969;
assign i[9727]= 16'he868;
assign i[9728]= 16'he7ba;
assign i[9729]= 16'he76a;
assign i[9730]= 16'he77e;
assign i[9731]= 16'he800;
assign i[9732]= 16'he8f4;
assign i[9733]= 16'hea60;
assign i[9734]= 16'hec43;
assign i[9735]= 16'hee9e;
assign i[9736]= 16'hf16b;
assign i[9737]= 16'hf4a5;
assign i[9738]= 16'hf841;
assign i[9739]= 16'hfc32;
assign i[9740]= 16'h65;
assign i[9741]= 16'h4cc;
assign i[9742]= 16'h94f;
assign i[9743]= 16'hdd8;
assign i[9744]= 16'h124f;
assign i[9745]= 16'h169d;
assign i[9746]= 16'h1aaa;
assign i[9747]= 16'h1e5f;
assign i[9748]= 16'h21a8;
assign i[9749]= 16'h2474;
assign i[9750]= 16'h26b5;
assign i[9751]= 16'h2860;
assign i[9752]= 16'h296f;
assign i[9753]= 16'h29e3;
assign i[9754]= 16'h29bd;
assign i[9755]= 16'h2908;
assign i[9756]= 16'h27d0;
assign i[9757]= 16'h2627;
assign i[9758]= 16'h2421;
assign i[9759]= 16'h21d7;
assign i[9760]= 16'h1f61;
assign i[9761]= 16'h1cdc;
assign i[9762]= 16'h1a61;
assign i[9763]= 16'h180c;
assign i[9764]= 16'h15f4;
assign i[9765]= 16'h142f;
assign i[9766]= 16'h12d1;
assign i[9767]= 16'h11e5;
assign i[9768]= 16'h1177;
assign i[9769]= 16'h118a;
assign i[9770]= 16'h121d;
assign i[9771]= 16'h132a;
assign i[9772]= 16'h14a6;
assign i[9773]= 16'h1682;
assign i[9774]= 16'h18aa;
assign i[9775]= 16'h1b08;
assign i[9776]= 16'h1d83;
assign i[9777]= 16'h2001;
assign i[9778]= 16'h2266;
assign i[9779]= 16'h249a;
assign i[9780]= 16'h2682;
assign i[9781]= 16'h280a;
assign i[9782]= 16'h291d;
assign i[9783]= 16'h29ac;
assign i[9784]= 16'h29ac;
assign i[9785]= 16'h2915;
assign i[9786]= 16'h27e7;
assign i[9787]= 16'h2622;
assign i[9788]= 16'h23cf;
assign i[9789]= 16'h20f8;
assign i[9790]= 16'h1dac;
assign i[9791]= 16'h19fd;
assign i[9792]= 16'h15fe;
assign i[9793]= 16'h11c6;
assign i[9794]= 16'hd6b;
assign i[9795]= 16'h905;
assign i[9796]= 16'h4a9;
assign i[9797]= 16'h6c;
assign i[9798]= 16'hfc64;
assign i[9799]= 16'hf89e;
assign i[9800]= 16'hf52c;
assign i[9801]= 16'hf218;
assign i[9802]= 16'hef6b;
assign i[9803]= 16'hed2c;
assign i[9804]= 16'heb5c;
assign i[9805]= 16'he9fd;
assign i[9806]= 16'he90b;
assign i[9807]= 16'he882;
assign i[9808]= 16'he85b;
assign i[9809]= 16'he88d;
assign i[9810]= 16'he910;
assign i[9811]= 16'he9d8;
assign i[9812]= 16'heada;
assign i[9813]= 16'hec0b;
assign i[9814]= 16'hed5e;
assign i[9815]= 16'heec8;
assign i[9816]= 16'hf03c;
assign i[9817]= 16'hf1b1;
assign i[9818]= 16'hf31a;
assign i[9819]= 16'hf46d;
assign i[9820]= 16'hf59f;
assign i[9821]= 16'hf6a8;
assign i[9822]= 16'hf77f;
assign i[9823]= 16'hf81c;
assign i[9824]= 16'hf876;
assign i[9825]= 16'hf889;
assign i[9826]= 16'hf850;
assign i[9827]= 16'hf7c5;
assign i[9828]= 16'hf6e8;
assign i[9829]= 16'hf5b8;
assign i[9830]= 16'hf437;
assign i[9831]= 16'hf268;
assign i[9832]= 16'hf051;
assign i[9833]= 16'hedfa;
assign i[9834]= 16'heb6e;
assign i[9835]= 16'he8ba;
assign i[9836]= 16'he5ed;
assign i[9837]= 16'he318;
assign i[9838]= 16'he04d;
assign i[9839]= 16'hdda0;
assign i[9840]= 16'hdb25;
assign i[9841]= 16'hd8f3;
assign i[9842]= 16'hd71c;
assign i[9843]= 16'hd5b6;
assign i[9844]= 16'hd4d1;
assign i[9845]= 16'hd47d;
assign i[9846]= 16'hd4c8;
assign i[9847]= 16'hd5bb;
assign i[9848]= 16'hd75c;
assign i[9849]= 16'hd9ac;
assign i[9850]= 16'hdcaa;
assign i[9851]= 16'he04d;
assign i[9852]= 16'he48c;
assign i[9853]= 16'he957;
assign i[9854]= 16'hee9b;
assign i[9855]= 16'hf442;
assign i[9856]= 16'hfa34;
assign i[9857]= 16'h54;
assign i[9858]= 16'h688;
assign i[9859]= 16'hcb4;
assign i[9860]= 16'h12bc;
assign i[9861]= 16'h1886;
assign i[9862]= 16'h1df9;
assign i[9863]= 16'h22ff;
assign i[9864]= 16'h2787;
assign i[9865]= 16'h2b82;
assign i[9866]= 16'h2ee6;
assign i[9867]= 16'h31ac;
assign i[9868]= 16'h33d4;
assign i[9869]= 16'h355f;
assign i[9870]= 16'h3654;
assign i[9871]= 16'h36bd;
assign i[9872]= 16'h36a7;
assign i[9873]= 16'h3621;
assign i[9874]= 16'h353b;
assign i[9875]= 16'h3408;
assign i[9876]= 16'h329a;
assign i[9877]= 16'h3101;
assign i[9878]= 16'h2f4e;
assign i[9879]= 16'h2d90;
assign i[9880]= 16'h2bd2;
assign i[9881]= 16'h2a1f;
assign i[9882]= 16'h287b;
assign i[9883]= 16'h26ec;
assign i[9884]= 16'h2572;
assign i[9885]= 16'h2409;
assign i[9886]= 16'h22af;
assign i[9887]= 16'h215a;
assign i[9888]= 16'h2003;
assign i[9889]= 16'h1ea0;
assign i[9890]= 16'h1d26;
assign i[9891]= 16'h1b8a;
assign i[9892]= 16'h19c1;
assign i[9893]= 16'h17c4;
assign i[9894]= 16'h158a;
assign i[9895]= 16'h130e;
assign i[9896]= 16'h104d;
assign i[9897]= 16'hd45;
assign i[9898]= 16'h9f9;
assign i[9899]= 16'h66d;
assign i[9900]= 16'h2a8;
assign i[9901]= 16'hfeb5;
assign i[9902]= 16'hfa9c;
assign i[9903]= 16'hf66c;
assign i[9904]= 16'hf232;
assign i[9905]= 16'hedfe;
assign i[9906]= 16'he9de;
assign i[9907]= 16'he5e2;
assign i[9908]= 16'he216;
assign i[9909]= 16'hde88;
assign i[9910]= 16'hdb43;
assign i[9911]= 16'hd850;
assign i[9912]= 16'hd5b6;
assign i[9913]= 16'hd37a;
assign i[9914]= 16'hd19f;
assign i[9915]= 16'hd024;
assign i[9916]= 16'hcf07;
assign i[9917]= 16'hce43;
assign i[9918]= 16'hcdd4;
assign i[9919]= 16'hcdb2;
assign i[9920]= 16'hcdd3;
assign i[9921]= 16'hce2f;
assign i[9922]= 16'hcebd;
assign i[9923]= 16'hcf72;
assign i[9924]= 16'hd046;
assign i[9925]= 16'hd130;
assign i[9926]= 16'hd229;
assign i[9927]= 16'hd32d;
assign i[9928]= 16'hd436;
assign i[9929]= 16'hd543;
assign i[9930]= 16'hd652;
assign i[9931]= 16'hd765;
assign i[9932]= 16'hd87e;
assign i[9933]= 16'hd9a2;
assign i[9934]= 16'hdad7;
assign i[9935]= 16'hdc21;
assign i[9936]= 16'hdd8a;
assign i[9937]= 16'hdf16;
assign i[9938]= 16'he0cf;
assign i[9939]= 16'he2bb;
assign i[9940]= 16'he4df;
assign i[9941]= 16'he740;
assign i[9942]= 16'he9e3;
assign i[9943]= 16'hecc7;
assign i[9944]= 16'hefee;
assign i[9945]= 16'hf355;
assign i[9946]= 16'hf6f6;
assign i[9947]= 16'hfacd;
assign i[9948]= 16'hfed0;
assign i[9949]= 16'h2f3;
assign i[9950]= 16'h72d;
assign i[9951]= 16'hb70;
assign i[9952]= 16'hfae;
assign i[9953]= 16'h13d7;
assign i[9954]= 16'h17dd;
assign i[9955]= 16'h1bb2;
assign i[9956]= 16'h1f49;
assign i[9957]= 16'h2295;
assign i[9958]= 16'h258c;
assign i[9959]= 16'h2827;
assign i[9960]= 16'h2a5f;
assign i[9961]= 16'h2c32;
assign i[9962]= 16'h2d9f;
assign i[9963]= 16'h2eaa;
assign i[9964]= 16'h2f57;
assign i[9965]= 16'h2faf;
assign i[9966]= 16'h2fbc;
assign i[9967]= 16'h2f8c;
assign i[9968]= 16'h2f2b;
assign i[9969]= 16'h2eaa;
assign i[9970]= 16'h2e17;
assign i[9971]= 16'h2d81;
assign i[9972]= 16'h2cf8;
assign i[9973]= 16'h2c87;
assign i[9974]= 16'h2c3b;
assign i[9975]= 16'h2c1a;
assign i[9976]= 16'h2c2c;
assign i[9977]= 16'h2c71;
assign i[9978]= 16'h2ce9;
assign i[9979]= 16'h2d8f;
assign i[9980]= 16'h2e5b;
assign i[9981]= 16'h2f41;
assign i[9982]= 16'h3033;
assign i[9983]= 16'h3120;
assign i[9984]= 16'h31f7;
assign i[9985]= 16'h32a3;
assign i[9986]= 16'h3313;
assign i[9987]= 16'h3333;
assign i[9988]= 16'h32f2;
assign i[9989]= 16'h3242;
assign i[9990]= 16'h3117;
assign i[9991]= 16'h2f69;
assign i[9992]= 16'h2d35;
assign i[9993]= 16'h2a7b;
assign i[9994]= 16'h2742;
assign i[9995]= 16'h2395;
assign i[9996]= 16'h1f83;
assign i[9997]= 16'h1b20;
assign i[9998]= 16'h1684;
assign i[9999]= 16'h11ca;
assign i[10000]= 16'hd0d;
assign i[10001]= 16'h86d;
assign i[10002]= 16'h407;
assign i[10003]= 16'hfff9;
assign i[10004]= 16'hfc5d;
assign i[10005]= 16'hf949;
assign i[10006]= 16'hf6d3;
assign i[10007]= 16'hf508;
assign i[10008]= 16'hf3f1;
assign i[10009]= 16'hf390;
assign i[10010]= 16'hf3e1;
assign i[10011]= 16'hf4d9;
assign i[10012]= 16'hf669;
assign i[10013]= 16'hf879;
assign i[10014]= 16'hfaef;
assign i[10015]= 16'hfdac;
assign i[10016]= 16'h8b;
assign i[10017]= 16'h36c;
assign i[10018]= 16'h628;
assign i[10019]= 16'h89e;
assign i[10020]= 16'haab;
assign i[10021]= 16'hc34;
assign i[10022]= 16'hd1e;
assign i[10023]= 16'hd59;
assign i[10024]= 16'hcd6;
assign i[10025]= 16'hb93;
assign i[10026]= 16'h990;
assign i[10027]= 16'h6d7;
assign i[10028]= 16'h379;
assign i[10029]= 16'hff8f;
assign i[10030]= 16'hfb34;
assign i[10031]= 16'hf68a;
assign i[10032]= 16'hf1b7;
assign i[10033]= 16'hece2;
assign i[10034]= 16'he833;
assign i[10035]= 16'he3d1;
assign i[10036]= 16'hdfe3;
assign i[10037]= 16'hdc89;
assign i[10038]= 16'hd9e0;
assign i[10039]= 16'hd7ff;
assign i[10040]= 16'hd6f6;
assign i[10041]= 16'hd6ce;
assign i[10042]= 16'hd789;
assign i[10043]= 16'hd920;
assign i[10044]= 16'hdb85;
assign i[10045]= 16'hdea4;
assign i[10046]= 16'he262;
assign i[10047]= 16'he6a0;
assign i[10048]= 16'heb3a;
assign i[10049]= 16'hf00b;
assign i[10050]= 16'hf4ea;
assign i[10051]= 16'hf9b2;
assign i[10052]= 16'hfe3d;
assign i[10053]= 16'h268;
assign i[10054]= 16'h616;
assign i[10055]= 16'h92e;
assign i[10056]= 16'hb9d;
assign i[10057]= 16'hd55;
assign i[10058]= 16'he51;
assign i[10059]= 16'he92;
assign i[10060]= 16'he1e;
assign i[10061]= 16'hd03;
assign i[10062]= 16'hb54;
assign i[10063]= 16'h928;
assign i[10064]= 16'h699;
assign i[10065]= 16'h3c5;
assign i[10066]= 16'hc7;
assign i[10067]= 16'hfdc0;
assign i[10068]= 16'hfaca;
assign i[10069]= 16'hf7ff;
assign i[10070]= 16'hf576;
assign i[10071]= 16'hf341;
assign i[10072]= 16'hf16e;
assign i[10073]= 16'hf004;
assign i[10074]= 16'hef08;
assign i[10075]= 16'hee76;
assign i[10076]= 16'hee47;
assign i[10077]= 16'hee6f;
assign i[10078]= 16'heedf;
assign i[10079]= 16'hef83;
assign i[10080]= 16'hf047;
assign i[10081]= 16'hf113;
assign i[10082]= 16'hf1d2;
assign i[10083]= 16'hf26f;
assign i[10084]= 16'hf2d4;
assign i[10085]= 16'hf2f2;
assign i[10086]= 16'hf2ba;
assign i[10087]= 16'hf223;
assign i[10088]= 16'hf127;
assign i[10089]= 16'hefc8;
assign i[10090]= 16'hee08;
assign i[10091]= 16'hebf3;
assign i[10092]= 16'he994;
assign i[10093]= 16'he6ff;
assign i[10094]= 16'he448;
assign i[10095]= 16'he187;
assign i[10096]= 16'hded6;
assign i[10097]= 16'hdc4e;
assign i[10098]= 16'hda0b;
assign i[10099]= 16'hd826;
assign i[10100]= 16'hd6b6;
assign i[10101]= 16'hd5d1;
assign i[10102]= 16'hd588;
assign i[10103]= 16'hd5e9;
assign i[10104]= 16'hd6fe;
assign i[10105]= 16'hd8cc;
assign i[10106]= 16'hdb53;
assign i[10107]= 16'hde8e;
assign i[10108]= 16'he274;
assign i[10109]= 16'he6f7;
assign i[10110]= 16'hec06;
assign i[10111]= 16'hf18c;
assign i[10112]= 16'hf772;
assign i[10113]= 16'hfd9d;
assign i[10114]= 16'h3f1;
assign i[10115]= 16'ha56;
assign i[10116]= 16'h10ae;
assign i[10117]= 16'h16de;
assign i[10118]= 16'h1cce;
assign i[10119]= 16'h2265;
assign i[10120]= 16'h278f;
assign i[10121]= 16'h2c3a;
assign i[10122]= 16'h3056;
assign i[10123]= 16'h33d7;
assign i[10124]= 16'h36b6;
assign i[10125]= 16'h38eb;
assign i[10126]= 16'h3a76;
assign i[10127]= 16'h3b56;
assign i[10128]= 16'h3b8f;
assign i[10129]= 16'h3b26;
assign i[10130]= 16'h3a23;
assign i[10131]= 16'h388f;
assign i[10132]= 16'h3673;
assign i[10133]= 16'h33db;
assign i[10134]= 16'h30d1;
assign i[10135]= 16'h2d62;
assign i[10136]= 16'h2997;
assign i[10137]= 16'h257d;
assign i[10138]= 16'h211d;
assign i[10139]= 16'h1c82;
assign i[10140]= 16'h17b4;
assign i[10141]= 16'h12bc;
assign i[10142]= 16'hda3;
assign i[10143]= 16'h86f;
assign i[10144]= 16'h32a;
assign i[10145]= 16'hfddc;
assign i[10146]= 16'hf88a;
assign i[10147]= 16'hf33f;
assign i[10148]= 16'hee02;
assign i[10149]= 16'he8de;
assign i[10150]= 16'he3dd;
assign i[10151]= 16'hdf0a;
assign i[10152]= 16'hda71;
assign i[10153]= 16'hd61e;
assign i[10154]= 16'hd21f;
assign i[10155]= 16'hce81;
assign i[10156]= 16'hcb51;
assign i[10157]= 16'hc89c;
assign i[10158]= 16'hc671;
assign i[10159]= 16'hc4d9;
assign i[10160]= 16'hc3e0;
assign i[10161]= 16'hc38e;
assign i[10162]= 16'hc3e9;
assign i[10163]= 16'hc4f6;
assign i[10164]= 16'hc6b6;
assign i[10165]= 16'hc926;
assign i[10166]= 16'hcc43;
assign i[10167]= 16'hd003;
assign i[10168]= 16'hd45a;
assign i[10169]= 16'hd93b;
assign i[10170]= 16'hde92;
assign i[10171]= 16'he44c;
assign i[10172]= 16'hea52;
assign i[10173]= 16'hf089;
assign i[10174]= 16'hf6d9;
assign i[10175]= 16'hfd26;
assign i[10176]= 16'h353;
assign i[10177]= 16'h946;
assign i[10178]= 16'hee6;
assign i[10179]= 16'h1419;
assign i[10180]= 16'h18c8;
assign i[10181]= 16'h1ce0;
assign i[10182]= 16'h2050;
assign i[10183]= 16'h230a;
assign i[10184]= 16'h2505;
assign i[10185]= 16'h263c;
assign i[10186]= 16'h26ac;
assign i[10187]= 16'h2657;
assign i[10188]= 16'h2543;
assign i[10189]= 16'h237b;
assign i[10190]= 16'h210a;
assign i[10191]= 16'h1e00;
assign i[10192]= 16'h1a6f;
assign i[10193]= 16'h166a;
assign i[10194]= 16'h1208;
assign i[10195]= 16'hd5e;
assign i[10196]= 16'h881;
assign i[10197]= 16'h389;
assign i[10198]= 16'hfe8b;
assign i[10199]= 16'hf99a;
assign i[10200]= 16'hf4ca;
assign i[10201]= 16'hf02b;
assign i[10202]= 16'hebcd;
assign i[10203]= 16'he7bc;
assign i[10204]= 16'he402;
assign i[10205]= 16'he0a8;
assign i[10206]= 16'hddb3;
assign i[10207]= 16'hdb27;
assign i[10208]= 16'hd906;
assign i[10209]= 16'hd74f;
assign i[10210]= 16'hd600;
assign i[10211]= 16'hd516;
assign i[10212]= 16'hd48b;
assign i[10213]= 16'hd45a;
assign i[10214]= 16'hd47d;
assign i[10215]= 16'hd4ec;
assign i[10216]= 16'hd5a0;
assign i[10217]= 16'hd691;
assign i[10218]= 16'hd7b7;
assign i[10219]= 16'hd90b;
assign i[10220]= 16'hda84;
assign i[10221]= 16'hdc1b;
assign i[10222]= 16'hddca;
assign i[10223]= 16'hdf88;
assign i[10224]= 16'he14f;
assign i[10225]= 16'he31a;
assign i[10226]= 16'he4e1;
assign i[10227]= 16'he6a1;
assign i[10228]= 16'he852;
assign i[10229]= 16'he9f2;
assign i[10230]= 16'heb7b;
assign i[10231]= 16'hece9;
assign i[10232]= 16'hee3a;
assign i[10233]= 16'hef6a;
assign i[10234]= 16'hf077;
assign i[10235]= 16'hf160;
assign i[10236]= 16'hf223;
assign i[10237]= 16'hf2bf;
assign i[10238]= 16'hf336;
assign i[10239]= 16'hf387;
assign i[10240]= 16'hf3b5;
assign i[10241]= 16'hf3c0;
assign i[10242]= 16'hf3ac;
assign i[10243]= 16'hf37b;
assign i[10244]= 16'hf330;
assign i[10245]= 16'hf2d0;
assign i[10246]= 16'hf25e;
assign i[10247]= 16'hf1df;
assign i[10248]= 16'hf157;
assign i[10249]= 16'hf0cb;
assign i[10250]= 16'hf040;
assign i[10251]= 16'hefb9;
assign i[10252]= 16'hef3d;
assign i[10253]= 16'heece;
assign i[10254]= 16'hee72;
assign i[10255]= 16'hee2d;
assign i[10256]= 16'hee02;
assign i[10257]= 16'hedf5;
assign i[10258]= 16'hee09;
assign i[10259]= 16'hee41;
assign i[10260]= 16'heea0;
assign i[10261]= 16'hef27;
assign i[10262]= 16'hefd8;
assign i[10263]= 16'hf0b4;
assign i[10264]= 16'hf1ba;
assign i[10265]= 16'hf2ea;
assign i[10266]= 16'hf442;
assign i[10267]= 16'hf5c1;
assign i[10268]= 16'hf763;
assign i[10269]= 16'hf924;
assign i[10270]= 16'hfb00;
assign i[10271]= 16'hfcf2;
assign i[10272]= 16'hfef2;
assign i[10273]= 16'hf9;
assign i[10274]= 16'h301;
assign i[10275]= 16'h503;
assign i[10276]= 16'h6f6;
assign i[10277]= 16'h8d3;
assign i[10278]= 16'ha92;
assign i[10279]= 16'hc2d;
assign i[10280]= 16'hd9d;
assign i[10281]= 16'hede;
assign i[10282]= 16'hfeb;
assign i[10283]= 16'h10c3;
assign i[10284]= 16'h1163;
assign i[10285]= 16'h11cd;
assign i[10286]= 16'h1201;
assign i[10287]= 16'h1203;
assign i[10288]= 16'h11d7;
assign i[10289]= 16'h1183;
assign i[10290]= 16'h110c;
assign i[10291]= 16'h1078;
assign i[10292]= 16'hfd0;
assign i[10293]= 16'hf18;
assign i[10294]= 16'he57;
assign i[10295]= 16'hd91;
assign i[10296]= 16'hccb;
assign i[10297]= 16'hc04;
assign i[10298]= 16'hb3f;
assign i[10299]= 16'ha79;
assign i[10300]= 16'h9af;
assign i[10301]= 16'h8da;
assign i[10302]= 16'h7f5;
assign i[10303]= 16'h6f7;
assign i[10304]= 16'h5d7;
assign i[10305]= 16'h48b;
assign i[10306]= 16'h309;
assign i[10307]= 16'h14a;
assign i[10308]= 16'hff46;
assign i[10309]= 16'hfcf7;
assign i[10310]= 16'hfa5a;
assign i[10311]= 16'hf770;
assign i[10312]= 16'hf43d;
assign i[10313]= 16'hf0c9;
assign i[10314]= 16'hed1f;
assign i[10315]= 16'he94e;
assign i[10316]= 16'he56a;
assign i[10317]= 16'he18a;
assign i[10318]= 16'hddc6;
assign i[10319]= 16'hda3b;
assign i[10320]= 16'hd705;
assign i[10321]= 16'hd440;
assign i[10322]= 16'hd20a;
assign i[10323]= 16'hd07b;
assign i[10324]= 16'hcfab;
assign i[10325]= 16'hcfad;
assign i[10326]= 16'hd08e;
assign i[10327]= 16'hd256;
assign i[10328]= 16'hd507;
assign i[10329]= 16'hd89b;
assign i[10330]= 16'hdd04;
assign i[10331]= 16'he22f;
assign i[10332]= 16'he801;
assign i[10333]= 16'hee59;
assign i[10334]= 16'hf511;
assign i[10335]= 16'hfbfd;
assign i[10336]= 16'h2f1;
assign i[10337]= 16'h9be;
assign i[10338]= 16'h1036;
assign i[10339]= 16'h162c;
assign i[10340]= 16'h1b77;
assign i[10341]= 16'h1ff2;
assign i[10342]= 16'h237f;
assign i[10343]= 16'h2607;
assign i[10344]= 16'h277d;
assign i[10345]= 16'h27da;
assign i[10346]= 16'h2724;
assign i[10347]= 16'h2567;
assign i[10348]= 16'h22ba;
assign i[10349]= 16'h1f3b;
assign i[10350]= 16'h1b11;
assign i[10351]= 16'h1667;
assign i[10352]= 16'h116e;
assign i[10353]= 16'hc58;
assign i[10354]= 16'h759;
assign i[10355]= 16'h2a3;
assign i[10356]= 16'hfe66;
assign i[10357]= 16'hfacb;
assign i[10358]= 16'hf7f8;
assign i[10359]= 16'hf608;
assign i[10360]= 16'hf50f;
assign i[10361]= 16'hf518;
assign i[10362]= 16'hf621;
assign i[10363]= 16'hf822;
assign i[10364]= 16'hfb06;
assign i[10365]= 16'hfeb0;
assign i[10366]= 16'h2fc;
assign i[10367]= 16'h7c0;
assign i[10368]= 16'hcca;
assign i[10369]= 16'h11e9;
assign i[10370]= 16'h16e8;
assign i[10371]= 16'h1b94;
assign i[10372]= 16'h1fbb;
assign i[10373]= 16'h2331;
assign i[10374]= 16'h25d1;
assign i[10375]= 16'h277b;
assign i[10376]= 16'h2819;
assign i[10377]= 16'h279d;
assign i[10378]= 16'h2605;
assign i[10379]= 16'h2357;
assign i[10380]= 16'h1fa2;
assign i[10381]= 16'h1afe;
assign i[10382]= 16'h158d;
assign i[10383]= 16'hf73;
assign i[10384]= 16'h8de;
assign i[10385]= 16'h1fa;
assign i[10386]= 16'hfafb;
assign i[10387]= 16'hf40e;
assign i[10388]= 16'hed63;
assign i[10389]= 16'he725;
assign i[10390]= 16'he17b;
assign i[10391]= 16'hdc85;
assign i[10392]= 16'hd85c;
assign i[10393]= 16'hd514;
assign i[10394]= 16'hd2b7;
assign i[10395]= 16'hd146;
assign i[10396]= 16'hd0bd;
assign i[10397]= 16'hd110;
assign i[10398]= 16'hd22c;
assign i[10399]= 16'hd3f9;
assign i[10400]= 16'hd65c;
assign i[10401]= 16'hd935;
assign i[10402]= 16'hdc64;
assign i[10403]= 16'hdfc8;
assign i[10404]= 16'he341;
assign i[10405]= 16'he6b0;
assign i[10406]= 16'he9fa;
assign i[10407]= 16'hed08;
assign i[10408]= 16'hefc6;
assign i[10409]= 16'hf226;
assign i[10410]= 16'hf41c;
assign i[10411]= 16'hf5a5;
assign i[10412]= 16'hf6c0;
assign i[10413]= 16'hf770;
assign i[10414]= 16'hf7bd;
assign i[10415]= 16'hf7b0;
assign i[10416]= 16'hf756;
assign i[10417]= 16'hf6be;
assign i[10418]= 16'hf5f6;
assign i[10419]= 16'hf50c;
assign i[10420]= 16'hf40f;
assign i[10421]= 16'hf30d;
assign i[10422]= 16'hf210;
assign i[10423]= 16'hf123;
assign i[10424]= 16'hf04e;
assign i[10425]= 16'hef95;
assign i[10426]= 16'heefc;
assign i[10427]= 16'hee86;
assign i[10428]= 16'hee32;
assign i[10429]= 16'hedff;
assign i[10430]= 16'hedea;
assign i[10431]= 16'hedef;
assign i[10432]= 16'hee0d;
assign i[10433]= 16'hee3d;
assign i[10434]= 16'hee7e;
assign i[10435]= 16'heecb;
assign i[10436]= 16'hef22;
assign i[10437]= 16'hef81;
assign i[10438]= 16'hefe4;
assign i[10439]= 16'hf04c;
assign i[10440]= 16'hf0b6;
assign i[10441]= 16'hf122;
assign i[10442]= 16'hf18e;
assign i[10443]= 16'hf1f8;
assign i[10444]= 16'hf260;
assign i[10445]= 16'hf2c3;
assign i[10446]= 16'hf31f;
assign i[10447]= 16'hf36f;
assign i[10448]= 16'hf3b1;
assign i[10449]= 16'hf3df;
assign i[10450]= 16'hf3f7;
assign i[10451]= 16'hf3f3;
assign i[10452]= 16'hf3d1;
assign i[10453]= 16'hf38c;
assign i[10454]= 16'hf324;
assign i[10455]= 16'hf297;
assign i[10456]= 16'hf1e8;
assign i[10457]= 16'hf118;
assign i[10458]= 16'hf02d;
assign i[10459]= 16'hef2e;
assign i[10460]= 16'hee25;
assign i[10461]= 16'hed1e;
assign i[10462]= 16'hec24;
assign i[10463]= 16'heb47;
assign i[10464]= 16'hea95;
assign i[10465]= 16'hea1f;
assign i[10466]= 16'he9f4;
assign i[10467]= 16'hea21;
assign i[10468]= 16'heab5;
assign i[10469]= 16'hebb8;
assign i[10470]= 16'hed33;
assign i[10471]= 16'hef2a;
assign i[10472]= 16'hf19e;
assign i[10473]= 16'hf48a;
assign i[10474]= 16'hf7e7;
assign i[10475]= 16'hfba9;
assign i[10476]= 16'hffbf;
assign i[10477]= 16'h416;
assign i[10478]= 16'h897;
assign i[10479]= 16'hd29;
assign i[10480]= 16'h11b1;
assign i[10481]= 16'h1613;
assign i[10482]= 16'h1a32;
assign i[10483]= 16'h1df3;
assign i[10484]= 16'h213e;
assign i[10485]= 16'h23fc;
assign i[10486]= 16'h261a;
assign i[10487]= 16'h278a;
assign i[10488]= 16'h2840;
assign i[10489]= 16'h2839;
assign i[10490]= 16'h2774;
assign i[10491]= 16'h25f7;
assign i[10492]= 16'h23cd;
assign i[10493]= 16'h2105;
assign i[10494]= 16'h1db2;
assign i[10495]= 16'h19eb;
assign i[10496]= 16'h15c8;
assign i[10497]= 16'h1167;
assign i[10498]= 16'hce2;
assign i[10499]= 16'h855;
assign i[10500]= 16'h3dc;
assign i[10501]= 16'hff91;
assign i[10502]= 16'hfb89;
assign i[10503]= 16'hf7d7;
assign i[10504]= 16'hf48b;
assign i[10505]= 16'hf1b2;
assign i[10506]= 16'hef53;
assign i[10507]= 16'hed6f;
assign i[10508]= 16'hec08;
assign i[10509]= 16'heb17;
assign i[10510]= 16'hea94;
assign i[10511]= 16'hea75;
assign i[10512]= 16'heaab;
assign i[10513]= 16'heb27;
assign i[10514]= 16'hebda;
assign i[10515]= 16'hecb2;
assign i[10516]= 16'heda1;
assign i[10517]= 16'hee96;
assign i[10518]= 16'hef86;
assign i[10519]= 16'hf063;
assign i[10520]= 16'hf125;
assign i[10521]= 16'hf1c4;
assign i[10522]= 16'hf23e;
assign i[10523]= 16'hf290;
assign i[10524]= 16'hf2bb;
assign i[10525]= 16'hf2c1;
assign i[10526]= 16'hf2a9;
assign i[10527]= 16'hf277;
assign i[10528]= 16'hf235;
assign i[10529]= 16'hf1ea;
assign i[10530]= 16'hf19f;
assign i[10531]= 16'hf15d;
assign i[10532]= 16'hf12d;
assign i[10533]= 16'hf117;
assign i[10534]= 16'hf121;
assign i[10535]= 16'hf152;
assign i[10536]= 16'hf1af;
assign i[10537]= 16'hf23a;
assign i[10538]= 16'hf2f6;
assign i[10539]= 16'hf3e5;
assign i[10540]= 16'hf505;
assign i[10541]= 16'hf657;
assign i[10542]= 16'hf7d7;
assign i[10543]= 16'hf984;
assign i[10544]= 16'hfb59;
assign i[10545]= 16'hfd54;
assign i[10546]= 16'hff70;
assign i[10547]= 16'h1a7;
assign i[10548]= 16'h3f8;
assign i[10549]= 16'h65d;
assign i[10550]= 16'h8d1;
assign i[10551]= 16'hb50;
assign i[10552]= 16'hdd5;
assign i[10553]= 16'h105d;
assign i[10554]= 16'h12e1;
assign i[10555]= 16'h155f;
assign i[10556]= 16'h17d0;
assign i[10557]= 16'h1a31;
assign i[10558]= 16'h1c7d;
assign i[10559]= 16'h1eaf;
assign i[10560]= 16'h20c3;
assign i[10561]= 16'h22b5;
assign i[10562]= 16'h2481;
assign i[10563]= 16'h2625;
assign i[10564]= 16'h279d;
assign i[10565]= 16'h28e8;
assign i[10566]= 16'h2a04;
assign i[10567]= 16'h2af2;
assign i[10568]= 16'h2bb2;
assign i[10569]= 16'h2c47;
assign i[10570]= 16'h2cb4;
assign i[10571]= 16'h2cfc;
assign i[10572]= 16'h2d24;
assign i[10573]= 16'h2d32;
assign i[10574]= 16'h2d2b;
assign i[10575]= 16'h2d17;
assign i[10576]= 16'h2cfb;
assign i[10577]= 16'h2cde;
assign i[10578]= 16'h2cc6;
assign i[10579]= 16'h2cb8;
assign i[10580]= 16'h2cb7;
assign i[10581]= 16'h2cc9;
assign i[10582]= 16'h2cee;
assign i[10583]= 16'h2d27;
assign i[10584]= 16'h2d73;
assign i[10585]= 16'h2dd1;
assign i[10586]= 16'h2e3c;
assign i[10587]= 16'h2eb0;
assign i[10588]= 16'h2f26;
assign i[10589]= 16'h2f98;
assign i[10590]= 16'h2ffe;
assign i[10591]= 16'h304f;
assign i[10592]= 16'h3083;
assign i[10593]= 16'h3092;
assign i[10594]= 16'h3074;
assign i[10595]= 16'h3021;
assign i[10596]= 16'h2f94;
assign i[10597]= 16'h2ec5;
assign i[10598]= 16'h2db2;
assign i[10599]= 16'h2c57;
assign i[10600]= 16'h2ab3;
assign i[10601]= 16'h28c5;
assign i[10602]= 16'h268e;
assign i[10603]= 16'h2411;
assign i[10604]= 16'h2152;
assign i[10605]= 16'h1e55;
assign i[10606]= 16'h1b20;
assign i[10607]= 16'h17bb;
assign i[10608]= 16'h142c;
assign i[10609]= 16'h107d;
assign i[10610]= 16'hcb5;
assign i[10611]= 16'h8de;
assign i[10612]= 16'h503;
assign i[10613]= 16'h12d;
assign i[10614]= 16'hfd68;
assign i[10615]= 16'hf9bc;
assign i[10616]= 16'hf636;
assign i[10617]= 16'hf2e1;
assign i[10618]= 16'hefc9;
assign i[10619]= 16'hecf8;
assign i[10620]= 16'hea79;
assign i[10621]= 16'he859;
assign i[10622]= 16'he6a0;
assign i[10623]= 16'he55a;
assign i[10624]= 16'he48e;
assign i[10625]= 16'he445;
assign i[10626]= 16'he484;
assign i[10627]= 16'he54f;
assign i[10628]= 16'he6a8;
assign i[10629]= 16'he88f;
assign i[10630]= 16'heaff;
assign i[10631]= 16'hedf2;
assign i[10632]= 16'hf15f;
assign i[10633]= 16'hf539;
assign i[10634]= 16'hf970;
assign i[10635]= 16'hfdf1;
assign i[10636]= 16'h2a6;
assign i[10637]= 16'h77a;
assign i[10638]= 16'hc51;
assign i[10639]= 16'h1110;
assign i[10640]= 16'h159e;
assign i[10641]= 16'h19de;
assign i[10642]= 16'h1db8;
assign i[10643]= 16'h2113;
assign i[10644]= 16'h23d9;
assign i[10645]= 16'h25f9;
assign i[10646]= 16'h2764;
assign i[10647]= 16'h2812;
assign i[10648]= 16'h27fe;
assign i[10649]= 16'h2728;
assign i[10650]= 16'h2598;
assign i[10651]= 16'h2359;
assign i[10652]= 16'h207c;
assign i[10653]= 16'h1d18;
assign i[10654]= 16'h1946;
assign i[10655]= 16'h1523;
assign i[10656]= 16'h10d0;
assign i[10657]= 16'hc6f;
assign i[10658]= 16'h822;
assign i[10659]= 16'h40a;
assign i[10660]= 16'h48;
assign i[10661]= 16'hfcfb;
assign i[10662]= 16'hfa3b;
assign i[10663]= 16'hf81f;
assign i[10664]= 16'hf6b8;
assign i[10665]= 16'hf613;
assign i[10666]= 16'hf633;
assign i[10667]= 16'hf71b;
assign i[10668]= 16'hf8c3;
assign i[10669]= 16'hfb21;
assign i[10670]= 16'hfe23;
assign i[10671]= 16'h1b5;
assign i[10672]= 16'h5c0;
assign i[10673]= 16'ha27;
assign i[10674]= 16'hecd;
assign i[10675]= 16'h1396;
assign i[10676]= 16'h1862;
assign i[10677]= 16'h1d16;
assign i[10678]= 16'h2197;
assign i[10679]= 16'h25cd;
assign i[10680]= 16'h29a3;
assign i[10681]= 16'h2d09;
assign i[10682]= 16'h2ff3;
assign i[10683]= 16'h3258;
assign i[10684]= 16'h3434;
assign i[10685]= 16'h3587;
assign i[10686]= 16'h3656;
assign i[10687]= 16'h36a9;
assign i[10688]= 16'h3688;
assign i[10689]= 16'h3601;
assign i[10690]= 16'h3521;
assign i[10691]= 16'h33f7;
assign i[10692]= 16'h3291;
assign i[10693]= 16'h30ff;
assign i[10694]= 16'h2f4e;
assign i[10695]= 16'h2d89;
assign i[10696]= 16'h2bbb;
assign i[10697]= 16'h29ec;
assign i[10698]= 16'h2822;
assign i[10699]= 16'h2661;
assign i[10700]= 16'h24ac;
assign i[10701]= 16'h2303;
assign i[10702]= 16'h2163;
assign i[10703]= 16'h1fcc;
assign i[10704]= 16'h1e39;
assign i[10705]= 16'h1ca6;
assign i[10706]= 16'h1b10;
assign i[10707]= 16'h1972;
assign i[10708]= 16'h17ca;
assign i[10709]= 16'h1616;
assign i[10710]= 16'h1453;
assign i[10711]= 16'h1281;
assign i[10712]= 16'h10a0;
assign i[10713]= 16'heb2;
assign i[10714]= 16'hcb9;
assign i[10715]= 16'hab9;
assign i[10716]= 16'h8b3;
assign i[10717]= 16'h6ad;
assign i[10718]= 16'h4a9;
assign i[10719]= 16'h2ac;
assign i[10720]= 16'hb8;
assign i[10721]= 16'hfed2;
assign i[10722]= 16'hfcf9;
assign i[10723]= 16'hfb30;
assign i[10724]= 16'hf979;
assign i[10725]= 16'hf7d5;
assign i[10726]= 16'hf642;
assign i[10727]= 16'hf4c3;
assign i[10728]= 16'hf356;
assign i[10729]= 16'hf1fe;
assign i[10730]= 16'hf0ba;
assign i[10731]= 16'hef8d;
assign i[10732]= 16'hee79;
assign i[10733]= 16'hed82;
assign i[10734]= 16'hecac;
assign i[10735]= 16'hebfd;
assign i[10736]= 16'heb79;
assign i[10737]= 16'heb27;
assign i[10738]= 16'heb0e;
assign i[10739]= 16'heb35;
assign i[10740]= 16'heba0;
assign i[10741]= 16'hec55;
assign i[10742]= 16'hed56;
assign i[10743]= 16'heea6;
assign i[10744]= 16'hf043;
assign i[10745]= 16'hf22a;
assign i[10746]= 16'hf455;
assign i[10747]= 16'hf6bb;
assign i[10748]= 16'hf951;
assign i[10749]= 16'hfc07;
assign i[10750]= 16'hfecf;
assign i[10751]= 16'h194;
assign i[10752]= 16'h444;
assign i[10753]= 16'h6ca;
assign i[10754]= 16'h913;
assign i[10755]= 16'hb09;
assign i[10756]= 16'hc9d;
assign i[10757]= 16'hdbe;
assign i[10758]= 16'he61;
assign i[10759]= 16'he7e;
assign i[10760]= 16'he12;
assign i[10761]= 16'hd1e;
assign i[10762]= 16'hba9;
assign i[10763]= 16'h9bf;
assign i[10764]= 16'h770;
assign i[10765]= 16'h4d1;
assign i[10766]= 16'h1fc;
assign i[10767]= 16'hff0e;
assign i[10768]= 16'hfc23;
assign i[10769]= 16'hf95c;
assign i[10770]= 16'hf6d7;
assign i[10771]= 16'hf4b4;
assign i[10772]= 16'hf30d;
assign i[10773]= 16'hf1fb;
assign i[10774]= 16'hf191;
assign i[10775]= 16'hf1dd;
assign i[10776]= 16'hf2e6;
assign i[10777]= 16'hf4ac;
assign i[10778]= 16'hf72a;
assign i[10779]= 16'hfa53;
assign i[10780]= 16'hfe12;
assign i[10781]= 16'h24c;
assign i[10782]= 16'h6e5;
assign i[10783]= 16'hbb7;
assign i[10784]= 16'h109d;
assign i[10785]= 16'h156f;
assign i[10786]= 16'h1a03;
assign i[10787]= 16'h1e35;
assign i[10788]= 16'h21df;
assign i[10789]= 16'h24e1;
assign i[10790]= 16'h2721;
assign i[10791]= 16'h288c;
assign i[10792]= 16'h2913;
assign i[10793]= 16'h28b3;
assign i[10794]= 16'h276e;
assign i[10795]= 16'h254f;
assign i[10796]= 16'h226a;
assign i[10797]= 16'h1ed7;
assign i[10798]= 16'h1ab8;
assign i[10799]= 16'h1631;
assign i[10800]= 16'h116c;
assign i[10801]= 16'hc92;
assign i[10802]= 16'h7d0;
assign i[10803]= 16'h351;
assign i[10804]= 16'hff3f;
assign i[10805]= 16'hfbbb;
assign i[10806]= 16'hf8e6;
assign i[10807]= 16'hf6da;
assign i[10808]= 16'hf5a9;
assign i[10809]= 16'hf55c;
assign i[10810]= 16'hf5f7;
assign i[10811]= 16'hf772;
assign i[10812]= 16'hf9c1;
assign i[10813]= 16'hfcce;
assign i[10814]= 16'h7d;
assign i[10815]= 16'h4af;
assign i[10816]= 16'h93f;
assign i[10817]= 16'he04;
assign i[10818]= 16'h12d5;
assign i[10819]= 16'h1788;
assign i[10820]= 16'h1bf6;
assign i[10821]= 16'h1ff9;
assign i[10822]= 16'h236f;
assign i[10823]= 16'h263d;
assign i[10824]= 16'h284b;
assign i[10825]= 16'h2989;
assign i[10826]= 16'h29ed;
assign i[10827]= 16'h2975;
assign i[10828]= 16'h2822;
assign i[10829]= 16'h2600;
assign i[10830]= 16'h231e;
assign i[10831]= 16'h1f8f;
assign i[10832]= 16'h1b6c;
assign i[10833]= 16'h16d1;
assign i[10834]= 16'h11db;
assign i[10835]= 16'hca7;
assign i[10836]= 16'h753;
assign i[10837]= 16'h1fd;
assign i[10838]= 16'hfcbf;
assign i[10839]= 16'hf7b0;
assign i[10840]= 16'hf2e5;
assign i[10841]= 16'hee6f;
assign i[10842]= 16'hea5b;
assign i[10843]= 16'he6b1;
assign i[10844]= 16'he376;
assign i[10845]= 16'he0aa;
assign i[10846]= 16'hde4c;
assign i[10847]= 16'hdc55;
assign i[10848]= 16'hdabf;
assign i[10849]= 16'hd97f;
assign i[10850]= 16'hd88b;
assign i[10851]= 16'hd7d9;
assign i[10852]= 16'hd75e;
assign i[10853]= 16'hd711;
assign i[10854]= 16'hd6e9;
assign i[10855]= 16'hd6e0;
assign i[10856]= 16'hd6f1;
assign i[10857]= 16'hd71a;
assign i[10858]= 16'hd75a;
assign i[10859]= 16'hd7b4;
assign i[10860]= 16'hd82a;
assign i[10861]= 16'hd8c3;
assign i[10862]= 16'hd985;
assign i[10863]= 16'hda77;
assign i[10864]= 16'hdba1;
assign i[10865]= 16'hdd0b;
assign i[10866]= 16'hdebc;
assign i[10867]= 16'he0b9;
assign i[10868]= 16'he307;
assign i[10869]= 16'he5a9;
assign i[10870]= 16'he89f;
assign i[10871]= 16'hebe8;
assign i[10872]= 16'hef7f;
assign i[10873]= 16'hf35c;
assign i[10874]= 16'hf777;
assign i[10875]= 16'hfbc5;
assign i[10876]= 16'h35;
assign i[10877]= 16'h4bc;
assign i[10878]= 16'h946;
assign i[10879]= 16'hdc3;
assign i[10880]= 16'h121f;
assign i[10881]= 16'h164b;
assign i[10882]= 16'h1a32;
assign i[10883]= 16'h1dc6;
assign i[10884]= 16'h20f8;
assign i[10885]= 16'h23ba;
assign i[10886]= 16'h2604;
assign i[10887]= 16'h27cc;
assign i[10888]= 16'h290e;
assign i[10889]= 16'h29c9;
assign i[10890]= 16'h29ff;
assign i[10891]= 16'h29b4;
assign i[10892]= 16'h28f1;
assign i[10893]= 16'h27c0;
assign i[10894]= 16'h262f;
assign i[10895]= 16'h244d;
assign i[10896]= 16'h222b;
assign i[10897]= 16'h1fdc;
assign i[10898]= 16'h1d72;
assign i[10899]= 16'h1b01;
assign i[10900]= 16'h189b;
assign i[10901]= 16'h1650;
assign i[10902]= 16'h1431;
assign i[10903]= 16'h124a;
assign i[10904]= 16'h10a7;
assign i[10905]= 16'hf4f;
assign i[10906]= 16'he46;
assign i[10907]= 16'hd8d;
assign i[10908]= 16'hd22;
assign i[10909]= 16'hcff;
assign i[10910]= 16'hd1b;
assign i[10911]= 16'hd6b;
assign i[10912]= 16'hde2;
assign i[10913]= 16'he6f;
assign i[10914]= 16'hf02;
assign i[10915]= 16'hf8b;
assign i[10916]= 16'hff9;
assign i[10917]= 16'h103c;
assign i[10918]= 16'h1046;
assign i[10919]= 16'h100c;
assign i[10920]= 16'hf84;
assign i[10921]= 16'hea9;
assign i[10922]= 16'hd79;
assign i[10923]= 16'hbf4;
assign i[10924]= 16'ha21;
assign i[10925]= 16'h809;
assign i[10926]= 16'h5b6;
assign i[10927]= 16'h338;
assign i[10928]= 16'ha0;
assign i[10929]= 16'hfe01;
assign i[10930]= 16'hfb6d;
assign i[10931]= 16'hf8f7;
assign i[10932]= 16'hf6b1;
assign i[10933]= 16'hf4ad;
assign i[10934]= 16'hf2f7;
assign i[10935]= 16'hf19a;
assign i[10936]= 16'hf09d;
assign i[10937]= 16'hf002;
assign i[10938]= 16'hefc8;
assign i[10939]= 16'hefe8;
assign i[10940]= 16'hf057;
assign i[10941]= 16'hf106;
assign i[10942]= 16'hf1e5;
assign i[10943]= 16'hf2de;
assign i[10944]= 16'hf3da;
assign i[10945]= 16'hf4c1;
assign i[10946]= 16'hf57e;
assign i[10947]= 16'hf5fa;
assign i[10948]= 16'hf620;
assign i[10949]= 16'hf5e1;
assign i[10950]= 16'hf531;
assign i[10951]= 16'hf407;
assign i[10952]= 16'hf263;
assign i[10953]= 16'hf047;
assign i[10954]= 16'hedbe;
assign i[10955]= 16'head7;
assign i[10956]= 16'he7a8;
assign i[10957]= 16'he448;
assign i[10958]= 16'he0d7;
assign i[10959]= 16'hdd74;
assign i[10960]= 16'hda41;
assign i[10961]= 16'hd761;
assign i[10962]= 16'hd4f5;
assign i[10963]= 16'hd31d;
assign i[10964]= 16'hd1f3;
assign i[10965]= 16'hd190;
assign i[10966]= 16'hd205;
assign i[10967]= 16'hd35b;
assign i[10968]= 16'hd598;
assign i[10969]= 16'hd8b7;
assign i[10970]= 16'hdcad;
assign i[10971]= 16'he168;
assign i[10972]= 16'he6ce;
assign i[10973]= 16'hecc0;
assign i[10974]= 16'hf31a;
assign i[10975]= 16'hf9b4;
assign i[10976]= 16'h63;
assign i[10977]= 16'h6fc;
assign i[10978]= 16'hd54;
assign i[10979]= 16'h1342;
assign i[10980]= 16'h189e;
assign i[10981]= 16'h1d48;
assign i[10982]= 16'h2123;
assign i[10983]= 16'h241a;
assign i[10984]= 16'h261f;
assign i[10985]= 16'h272a;
assign i[10986]= 16'h273c;
assign i[10987]= 16'h265c;
assign i[10988]= 16'h249c;
assign i[10989]= 16'h220e;
assign i[10990]= 16'h1ed0;
assign i[10991]= 16'h1b01;
assign i[10992]= 16'h16c3;
assign i[10993]= 16'h123c;
assign i[10994]= 16'hd92;
assign i[10995]= 16'h8ea;
assign i[10996]= 16'h469;
assign i[10997]= 16'h2f;
assign i[10998]= 16'hfc5c;
assign i[10999]= 16'hf907;
assign i[11000]= 16'hf644;
assign i[11001]= 16'hf421;
assign i[11002]= 16'hf2a8;
assign i[11003]= 16'hf1db;
assign i[11004]= 16'hf1b8;
assign i[11005]= 16'hf236;
assign i[11006]= 16'hf349;
assign i[11007]= 16'hf4df;
assign i[11008]= 16'hf6e6;
assign i[11009]= 16'hf946;
assign i[11010]= 16'hfbe6;
assign i[11011]= 16'hfeae;
assign i[11012]= 16'h182;
assign i[11013]= 16'h44b;
assign i[11014]= 16'h6f1;
assign i[11015]= 16'h95e;
assign i[11016]= 16'hb7f;
assign i[11017]= 16'hd41;
assign i[11018]= 16'he98;
assign i[11019]= 16'hf78;
assign i[11020]= 16'hfdb;
assign i[11021]= 16'hfba;
assign i[11022]= 16'hf16;
assign i[11023]= 16'hdef;
assign i[11024]= 16'hc49;
assign i[11025]= 16'ha2c;
assign i[11026]= 16'h7a1;
assign i[11027]= 16'h4b3;
assign i[11028]= 16'h16e;
assign i[11029]= 16'hfde2;
assign i[11030]= 16'hfa1c;
assign i[11031]= 16'hf62e;
assign i[11032]= 16'hf229;
assign i[11033]= 16'hee1e;
assign i[11034]= 16'hea20;
assign i[11035]= 16'he640;
assign i[11036]= 16'he290;
assign i[11037]= 16'hdf21;
assign i[11038]= 16'hdc03;
assign i[11039]= 16'hd946;
assign i[11040]= 16'hd6f7;
assign i[11041]= 16'hd523;
assign i[11042]= 16'hd3d5;
assign i[11043]= 16'hd315;
assign i[11044]= 16'hd2ea;
assign i[11045]= 16'hd359;
assign i[11046]= 16'hd464;
assign i[11047]= 16'hd60a;
assign i[11048]= 16'hd847;
assign i[11049]= 16'hdb17;
assign i[11050]= 16'hde70;
assign i[11051]= 16'he24a;
assign i[11052]= 16'he697;
assign i[11053]= 16'heb49;
assign i[11054]= 16'hf050;
assign i[11055]= 16'hf59b;
assign i[11056]= 16'hfb18;
assign i[11057]= 16'hb4;
assign i[11058]= 16'h65e;
assign i[11059]= 16'hc02;
assign i[11060]= 16'h118e;
assign i[11061]= 16'h16f0;
assign i[11062]= 16'h1c19;
assign i[11063]= 16'h20f9;
assign i[11064]= 16'h2584;
assign i[11065]= 16'h29ab;
assign i[11066]= 16'h2d66;
assign i[11067]= 16'h30ac;
assign i[11068]= 16'h3376;
assign i[11069]= 16'h35bf;
assign i[11070]= 16'h3783;
assign i[11071]= 16'h38c0;
assign i[11072]= 16'h3978;
assign i[11073]= 16'h39ac;
assign i[11074]= 16'h395e;
assign i[11075]= 16'h3895;
assign i[11076]= 16'h3756;
assign i[11077]= 16'h35aa;
assign i[11078]= 16'h339c;
assign i[11079]= 16'h3136;
assign i[11080]= 16'h2e85;
assign i[11081]= 16'h2b98;
assign i[11082]= 16'h287e;
assign i[11083]= 16'h2549;
assign i[11084]= 16'h220a;
assign i[11085]= 16'h1ed5;
assign i[11086]= 16'h1bbb;
assign i[11087]= 16'h18d0;
assign i[11088]= 16'h1626;
assign i[11089]= 16'h13cf;
assign i[11090]= 16'h11da;
assign i[11091]= 16'h1055;
assign i[11092]= 16'hf4c;
assign i[11093]= 16'hec5;
assign i[11094]= 16'hec6;
assign i[11095]= 16'hf4f;
assign i[11096]= 16'h105d;
assign i[11097]= 16'h11e8;
assign i[11098]= 16'h13e3;
assign i[11099]= 16'h163e;
assign i[11100]= 16'h18e5;
assign i[11101]= 16'h1bc0;
assign i[11102]= 16'h1eb5;
assign i[11103]= 16'h21a8;
assign i[11104]= 16'h247c;
assign i[11105]= 16'h2714;
assign i[11106]= 16'h2952;
assign i[11107]= 16'h2b1d;
assign i[11108]= 16'h2c5f;
assign i[11109]= 16'h2d02;
assign i[11110]= 16'h2cfa;
assign i[11111]= 16'h2c3d;
assign i[11112]= 16'h2ac8;
assign i[11113]= 16'h28a0;
assign i[11114]= 16'h25cd;
assign i[11115]= 16'h2262;
assign i[11116]= 16'h1e73;
assign i[11117]= 16'h1a1c;
assign i[11118]= 16'h157d;
assign i[11119]= 16'h10b9;
assign i[11120]= 16'hbf6;
assign i[11121]= 16'h759;
assign i[11122]= 16'h308;
assign i[11123]= 16'hff28;
assign i[11124]= 16'hfbd8;
assign i[11125]= 16'hf933;
assign i[11126]= 16'hf751;
assign i[11127]= 16'hf642;
assign i[11128]= 16'hf60d;
assign i[11129]= 16'hf6b6;
assign i[11130]= 16'hf835;
assign i[11131]= 16'hfa7d;
assign i[11132]= 16'hfd78;
assign i[11133]= 16'h10c;
assign i[11134]= 16'h518;
assign i[11135]= 16'h978;
assign i[11136]= 16'he02;
assign i[11137]= 16'h128f;
assign i[11138]= 16'h16f3;
assign i[11139]= 16'h1b05;
assign i[11140]= 16'h1ea0;
assign i[11141]= 16'h21a1;
assign i[11142]= 16'h23ea;
assign i[11143]= 16'h2563;
assign i[11144]= 16'h25fa;
assign i[11145]= 16'h25a5;
assign i[11146]= 16'h2460;
assign i[11147]= 16'h222e;
assign i[11148]= 16'h1f1a;
assign i[11149]= 16'h1b33;
assign i[11150]= 16'h1691;
assign i[11151]= 16'h114e;
assign i[11152]= 16'hb87;
assign i[11153]= 16'h560;
assign i[11154]= 16'hfefc;
assign i[11155]= 16'hf87c;
assign i[11156]= 16'hf206;
assign i[11157]= 16'hebbc;
assign i[11158]= 16'he5bf;
assign i[11159]= 16'he02c;
assign i[11160]= 16'hdb1f;
assign i[11161]= 16'hd6af;
assign i[11162]= 16'hd2ef;
assign i[11163]= 16'hcfef;
assign i[11164]= 16'hcdbb;
assign i[11165]= 16'hcc59;
assign i[11166]= 16'hcbcf;
assign i[11167]= 16'hcc1b;
assign i[11168]= 16'hcd3b;
assign i[11169]= 16'hcf2a;
assign i[11170]= 16'hd1dd;
assign i[11171]= 16'hd548;
assign i[11172]= 16'hd95f;
assign i[11173]= 16'hde0e;
assign i[11174]= 16'he345;
assign i[11175]= 16'he8ed;
assign i[11176]= 16'heef0;
assign i[11177]= 16'hf534;
assign i[11178]= 16'hfb9e;
assign i[11179]= 16'h212;
assign i[11180]= 16'h874;
assign i[11181]= 16'hea5;
assign i[11182]= 16'h1486;
assign i[11183]= 16'h19f8;
assign i[11184]= 16'h1ede;
assign i[11185]= 16'h231c;
assign i[11186]= 16'h2698;
assign i[11187]= 16'h293a;
assign i[11188]= 16'h2af0;
assign i[11189]= 16'h2bac;
assign i[11190]= 16'h2b65;
assign i[11191]= 16'h2a17;
assign i[11192]= 16'h27c7;
assign i[11193]= 16'h247f;
assign i[11194]= 16'h2052;
assign i[11195]= 16'h1b56;
assign i[11196]= 16'h15ac;
assign i[11197]= 16'hf79;
assign i[11198]= 16'h8e6;
assign i[11199]= 16'h221;
assign i[11200]= 16'hfb5d;
assign i[11201]= 16'hf4c9;
assign i[11202]= 16'hee99;
assign i[11203]= 16'he8fc;
assign i[11204]= 16'he41f;
assign i[11205]= 16'he029;
assign i[11206]= 16'hdd3b;
assign i[11207]= 16'hdb6f;
assign i[11208]= 16'hdad4;
assign i[11209]= 16'hdb71;
assign i[11210]= 16'hdd42;
assign i[11211]= 16'he03b;
assign i[11212]= 16'he443;
assign i[11213]= 16'he93b;
assign i[11214]= 16'heef8;
assign i[11215]= 16'hf54b;
assign i[11216]= 16'hfc00;
assign i[11217]= 16'h2db;
assign i[11218]= 16'h9a4;
assign i[11219]= 16'h1020;
assign i[11220]= 16'h1617;
assign i[11221]= 16'h1b54;
assign i[11222]= 16'h1fab;
assign i[11223]= 16'h22f4;
assign i[11224]= 16'h2513;
assign i[11225]= 16'h25f4;
assign i[11226]= 16'h258f;
assign i[11227]= 16'h23e6;
assign i[11228]= 16'h2107;
assign i[11229]= 16'h1d08;
assign i[11230]= 16'h180a;
assign i[11231]= 16'h1235;
assign i[11232]= 16'hbba;
assign i[11233]= 16'h4cd;
assign i[11234]= 16'hfda5;
assign i[11235]= 16'hf67a;
assign i[11236]= 16'hef85;
assign i[11237]= 16'he8fb;
assign i[11238]= 16'he30d;
assign i[11239]= 16'hdde7;
assign i[11240]= 16'hd9ab;
assign i[11241]= 16'hd677;
assign i[11242]= 16'hd45e;
assign i[11243]= 16'hd369;
assign i[11244]= 16'hd39a;
assign i[11245]= 16'hd4e9;
assign i[11246]= 16'hd747;
assign i[11247]= 16'hda9c;
assign i[11248]= 16'hdecb;
assign i[11249]= 16'he3b2;
assign i[11250]= 16'he92d;
assign i[11251]= 16'hef13;
assign i[11252]= 16'hf53d;
assign i[11253]= 16'hfb83;
assign i[11254]= 16'h1c0;
assign i[11255]= 16'h7d3;
assign i[11256]= 16'hd9e;
assign i[11257]= 16'h1306;
assign i[11258]= 16'h17f7;
assign i[11259]= 16'h1c61;
assign i[11260]= 16'h203c;
assign i[11261]= 16'h2380;
assign i[11262]= 16'h262f;
assign i[11263]= 16'h2849;
assign i[11264]= 16'h29d8;
assign i[11265]= 16'h2ae2;
assign i[11266]= 16'h2b73;
assign i[11267]= 16'h2b96;
assign i[11268]= 16'h2b56;
assign i[11269]= 16'h2ac0;
assign i[11270]= 16'h29dc;
assign i[11271]= 16'h28b4;
assign i[11272]= 16'h274f;
assign i[11273]= 16'h25b2;
assign i[11274]= 16'h23df;
assign i[11275]= 16'h21da;
assign i[11276]= 16'h1fa1;
assign i[11277]= 16'h1d36;
assign i[11278]= 16'h1a95;
assign i[11279]= 16'h17be;
assign i[11280]= 16'h14af;
assign i[11281]= 16'h1169;
assign i[11282]= 16'hded;
assign i[11283]= 16'ha3c;
assign i[11284]= 16'h65c;
assign i[11285]= 16'h253;
assign i[11286]= 16'hfe2b;
assign i[11287]= 16'hf9eb;
assign i[11288]= 16'hf5a1;
assign i[11289]= 16'hf15c;
assign i[11290]= 16'hed29;
assign i[11291]= 16'he918;
assign i[11292]= 16'he539;
assign i[11293]= 16'he19d;
assign i[11294]= 16'hde52;
assign i[11295]= 16'hdb65;
assign i[11296]= 16'hd8e3;
assign i[11297]= 16'hd6d6;
assign i[11298]= 16'hd545;
assign i[11299]= 16'hd437;
assign i[11300]= 16'hd3ad;
assign i[11301]= 16'hd3a8;
assign i[11302]= 16'hd426;
assign i[11303]= 16'hd521;
assign i[11304]= 16'hd693;
assign i[11305]= 16'hd873;
assign i[11306]= 16'hdab6;
assign i[11307]= 16'hdd52;
assign i[11308]= 16'he039;
assign i[11309]= 16'he360;
assign i[11310]= 16'he6b9;
assign i[11311]= 16'hea38;
assign i[11312]= 16'hedd1;
assign i[11313]= 16'hf178;
assign i[11314]= 16'hf522;
assign i[11315]= 16'hf8c6;
assign i[11316]= 16'hfc59;
assign i[11317]= 16'hffd4;
assign i[11318]= 16'h32e;
assign i[11319]= 16'h662;
assign i[11320]= 16'h967;
assign i[11321]= 16'hc37;
assign i[11322]= 16'hecd;
assign i[11323]= 16'h1121;
assign i[11324]= 16'h132f;
assign i[11325]= 16'h14f0;
assign i[11326]= 16'h165e;
assign i[11327]= 16'h1775;
assign i[11328]= 16'h182f;
assign i[11329]= 16'h1889;
assign i[11330]= 16'h187f;
assign i[11331]= 16'h180f;
assign i[11332]= 16'h1739;
assign i[11333]= 16'h15ff;
assign i[11334]= 16'h1464;
assign i[11335]= 16'h126d;
assign i[11336]= 16'h1022;
assign i[11337]= 16'hd8f;
assign i[11338]= 16'hac0;
assign i[11339]= 16'h7c4;
assign i[11340]= 16'h4ad;
assign i[11341]= 16'h18f;
assign i[11342]= 16'hfe7d;
assign i[11343]= 16'hfb8d;
assign i[11344]= 16'hf8d5;
assign i[11345]= 16'hf669;
assign i[11346]= 16'hf45f;
assign i[11347]= 16'hf2ca;
assign i[11348]= 16'hf1b8;
assign i[11349]= 16'hf138;
assign i[11350]= 16'hf153;
assign i[11351]= 16'hf20f;
assign i[11352]= 16'hf36d;
assign i[11353]= 16'hf569;
assign i[11354]= 16'hf7fb;
assign i[11355]= 16'hfb16;
assign i[11356]= 16'hfea9;
assign i[11357]= 16'h29e;
assign i[11358]= 16'h6de;
assign i[11359]= 16'hb4e;
assign i[11360]= 16'hfd0;
assign i[11361]= 16'h1447;
assign i[11362]= 16'h1894;
assign i[11363]= 16'h1c9b;
assign i[11364]= 16'h2042;
assign i[11365]= 16'h2370;
assign i[11366]= 16'h2613;
assign i[11367]= 16'h2819;
assign i[11368]= 16'h297b;
assign i[11369]= 16'h2a32;
assign i[11370]= 16'h2a41;
assign i[11371]= 16'h29af;
assign i[11372]= 16'h2887;
assign i[11373]= 16'h26dc;
assign i[11374]= 16'h24c5;
assign i[11375]= 16'h225a;
assign i[11376]= 16'h1fba;
assign i[11377]= 16'h1d03;
assign i[11378]= 16'h1a53;
assign i[11379]= 16'h17cb;
assign i[11380]= 16'h1586;
assign i[11381]= 16'h139e;
assign i[11382]= 16'h122a;
assign i[11383]= 16'h113b;
assign i[11384]= 16'h10dc;
assign i[11385]= 16'h1113;
assign i[11386]= 16'h11df;
assign i[11387]= 16'h1338;
assign i[11388]= 16'h1510;
assign i[11389]= 16'h1755;
assign i[11390]= 16'h19ec;
assign i[11391]= 16'h1cba;
assign i[11392]= 16'h1f9c;
assign i[11393]= 16'h2272;
assign i[11394]= 16'h2516;
assign i[11395]= 16'h2766;
assign i[11396]= 16'h2941;
assign i[11397]= 16'h2a88;
assign i[11398]= 16'h2b22;
assign i[11399]= 16'h2af8;
assign i[11400]= 16'h29fd;
assign i[11401]= 16'h2827;
assign i[11402]= 16'h2577;
assign i[11403]= 16'h21f1;
assign i[11404]= 16'h1da3;
assign i[11405]= 16'h18a0;
assign i[11406]= 16'h1301;
assign i[11407]= 16'hce4;
assign i[11408]= 16'h66c;
assign i[11409]= 16'hffbe;
assign i[11410]= 16'hf8fe;
assign i[11411]= 16'hf255;
assign i[11412]= 16'hebe5;
assign i[11413]= 16'he5d3;
assign i[11414]= 16'he03b;
assign i[11415]= 16'hdb39;
assign i[11416]= 16'hd6de;
assign i[11417]= 16'hd33a;
assign i[11418]= 16'hd053;
assign i[11419]= 16'hce29;
assign i[11420]= 16'hccb7;
assign i[11421]= 16'hcbef;
assign i[11422]= 16'hcbc0;
assign i[11423]= 16'hcc14;
assign i[11424]= 16'hccd0;
assign i[11425]= 16'hcdd9;
assign i[11426]= 16'hcf12;
assign i[11427]= 16'hd05c;
assign i[11428]= 16'hd19e;
assign i[11429]= 16'hd2be;
assign i[11430]= 16'hd3a6;
assign i[11431]= 16'hd447;
assign i[11432]= 16'hd496;
assign i[11433]= 16'hd48c;
assign i[11434]= 16'hd42b;
assign i[11435]= 16'hd37a;
assign i[11436]= 16'hd284;
assign i[11437]= 16'hd15b;
assign i[11438]= 16'hd016;
assign i[11439]= 16'hcecc;
assign i[11440]= 16'hcd9b;
assign i[11441]= 16'hcc9e;
assign i[11442]= 16'hcbf3;
assign i[11443]= 16'hcbb4;
assign i[11444]= 16'hcbfb;
assign i[11445]= 16'hccdd;
assign i[11446]= 16'hce69;
assign i[11447]= 16'hd0ac;
assign i[11448]= 16'hd3a9;
assign i[11449]= 16'hd760;
assign i[11450]= 16'hdbc9;
assign i[11451]= 16'he0d5;
assign i[11452]= 16'he66f;
assign i[11453]= 16'hec7d;
assign i[11454]= 16'hf2e1;
assign i[11455]= 16'hf979;
assign i[11456]= 16'h1f;
assign i[11457]= 16'h6ad;
assign i[11458]= 16'hcfe;
assign i[11459]= 16'h12eb;
assign i[11460]= 16'h1852;
assign i[11461]= 16'h1d13;
assign i[11462]= 16'h2113;
assign i[11463]= 16'h243d;
assign i[11464]= 16'h2681;
assign i[11465]= 16'h27d5;
assign i[11466]= 16'h2838;
assign i[11467]= 16'h27ac;
assign i[11468]= 16'h263d;
assign i[11469]= 16'h23fa;
assign i[11470]= 16'h20f9;
assign i[11471]= 16'h1d54;
assign i[11472]= 16'h1929;
assign i[11473]= 16'h1498;
assign i[11474]= 16'hfc3;
assign i[11475]= 16'hacb;
assign i[11476]= 16'h5d3;
assign i[11477]= 16'hf9;
assign i[11478]= 16'hfc5d;
assign i[11479]= 16'hf815;
assign i[11480]= 16'hf439;
assign i[11481]= 16'hf0d8;
assign i[11482]= 16'hee01;
assign i[11483]= 16'hebba;
assign i[11484]= 16'hea04;
assign i[11485]= 16'he8df;
assign i[11486]= 16'he843;
assign i[11487]= 16'he827;
assign i[11488]= 16'he87c;
assign i[11489]= 16'he933;
assign i[11490]= 16'hea3b;
assign i[11491]= 16'heb82;
assign i[11492]= 16'hecf5;
assign i[11493]= 16'hee85;
assign i[11494]= 16'hf021;
assign i[11495]= 16'hf1bc;
assign i[11496]= 16'hf34b;
assign i[11497]= 16'hf4c7;
assign i[11498]= 16'hf62b;
assign i[11499]= 16'hf775;
assign i[11500]= 16'hf8a9;
assign i[11501]= 16'hf9ca;
assign i[11502]= 16'hfae0;
assign i[11503]= 16'hfbf5;
assign i[11504]= 16'hfd12;
assign i[11505]= 16'hfe45;
assign i[11506]= 16'hff98;
assign i[11507]= 16'h115;
assign i[11508]= 16'h2c8;
assign i[11509]= 16'h4b9;
assign i[11510]= 16'h6eb;
assign i[11511]= 16'h960;
assign i[11512]= 16'hc19;
assign i[11513]= 16'hf0e;
assign i[11514]= 16'h1238;
assign i[11515]= 16'h1589;
assign i[11516]= 16'h18f2;
assign i[11517]= 16'h1c60;
assign i[11518]= 16'h1fbd;
assign i[11519]= 16'h22f1;
assign i[11520]= 16'h25e5;
assign i[11521]= 16'h2880;
assign i[11522]= 16'h2aa9;
assign i[11523]= 16'h2c4a;
assign i[11524]= 16'h2d4f;
assign i[11525]= 16'h2da6;
assign i[11526]= 16'h2d43;
assign i[11527]= 16'h2c1c;
assign i[11528]= 16'h2a2e;
assign i[11529]= 16'h277a;
assign i[11530]= 16'h2407;
assign i[11531]= 16'h1fe0;
assign i[11532]= 16'h1b18;
assign i[11533]= 16'h15c2;
assign i[11534]= 16'hff9;
assign i[11535]= 16'h9da;
assign i[11536]= 16'h383;
assign i[11537]= 16'hfd16;
assign i[11538]= 16'hf6b1;
assign i[11539]= 16'hf075;
assign i[11540]= 16'hea81;
assign i[11541]= 16'he4ef;
assign i[11542]= 16'hdfd9;
assign i[11543]= 16'hdb50;
assign i[11544]= 16'hd764;
assign i[11545]= 16'hd41e;
assign i[11546]= 16'hd182;
assign i[11547]= 16'hcf8e;
assign i[11548]= 16'hce3a;
assign i[11549]= 16'hcd7b;
assign i[11550]= 16'hcd3f;
assign i[11551]= 16'hcd73;
assign i[11552]= 16'hce01;
assign i[11553]= 16'hcecf;
assign i[11554]= 16'hcfc4;
assign i[11555]= 16'hd0c9;
assign i[11556]= 16'hd1c4;
assign i[11557]= 16'hd2a2;
assign i[11558]= 16'hd352;
assign i[11559]= 16'hd3c4;
assign i[11560]= 16'hd3f1;
assign i[11561]= 16'hd3d5;
assign i[11562]= 16'hd371;
assign i[11563]= 16'hd2ca;
assign i[11564]= 16'hd1ed;
assign i[11565]= 16'hd0e9;
assign i[11566]= 16'hcfd0;
assign i[11567]= 16'hceb9;
assign i[11568]= 16'hcdbd;
assign i[11569]= 16'hccf3;
assign i[11570]= 16'hcc76;
assign i[11571]= 16'hcc5e;
assign i[11572]= 16'hccbf;
assign i[11573]= 16'hcdac;
assign i[11574]= 16'hcf34;
assign i[11575]= 16'hd162;
assign i[11576]= 16'hd439;
assign i[11577]= 16'hd7b9;
assign i[11578]= 16'hdbdb;
assign i[11579]= 16'he095;
assign i[11580]= 16'he5d5;
assign i[11581]= 16'heb86;
assign i[11582]= 16'hf18e;
assign i[11583]= 16'hf7d0;
assign i[11584]= 16'hfe2f;
assign i[11585]= 16'h488;
assign i[11586]= 16'habe;
assign i[11587]= 16'h10b1;
assign i[11588]= 16'h1643;
assign i[11589]= 16'h1b5a;
assign i[11590]= 16'h1fdf;
assign i[11591]= 16'h23bf;
assign i[11592]= 16'h26ec;
assign i[11593]= 16'h295d;
assign i[11594]= 16'h2b0f;
assign i[11595]= 16'h2c04;
assign i[11596]= 16'h2c41;
assign i[11597]= 16'h2bd2;
assign i[11598]= 16'h2ac6;
assign i[11599]= 16'h292f;
assign i[11600]= 16'h2724;
assign i[11601]= 16'h24ba;
assign i[11602]= 16'h220b;
assign i[11603]= 16'h1f2e;
assign i[11604]= 16'h1c3c;
assign i[11605]= 16'h194c;
assign i[11606]= 16'h1672;
assign i[11607]= 16'h13c1;
assign i[11608]= 16'h1149;
assign i[11609]= 16'hf17;
assign i[11610]= 16'hd34;
assign i[11611]= 16'hba7;
assign i[11612]= 16'ha72;
assign i[11613]= 16'h995;
assign i[11614]= 16'h90e;
assign i[11615]= 16'h8d7;
assign i[11616]= 16'h8ea;
assign i[11617]= 16'h93d;
assign i[11618]= 16'h9c6;
assign i[11619]= 16'ha7b;
assign i[11620]= 16'hb50;
assign i[11621]= 16'hc3b;
assign i[11622]= 16'hd31;
assign i[11623]= 16'he29;
assign i[11624]= 16'hf19;
assign i[11625]= 16'hff9;
assign i[11626]= 16'h10c3;
assign i[11627]= 16'h1172;
assign i[11628]= 16'h1201;
assign i[11629]= 16'h126d;
assign i[11630]= 16'h12b6;
assign i[11631]= 16'h12da;
assign i[11632]= 16'h12da;
assign i[11633]= 16'h12b7;
assign i[11634]= 16'h1273;
assign i[11635]= 16'h1211;
assign i[11636]= 16'h1196;
assign i[11637]= 16'h1104;
assign i[11638]= 16'h1060;
assign i[11639]= 16'hfaf;
assign i[11640]= 16'hef7;
assign i[11641]= 16'he3d;
assign i[11642]= 16'hd86;
assign i[11643]= 16'hcd9;
assign i[11644]= 16'hc3b;
assign i[11645]= 16'hbb3;
assign i[11646]= 16'hb46;
assign i[11647]= 16'hafa;
assign i[11648]= 16'had4;
assign i[11649]= 16'had9;
assign i[11650]= 16'hb0c;
assign i[11651]= 16'hb71;
assign i[11652]= 16'hc0b;
assign i[11653]= 16'hcda;
assign i[11654]= 16'hddf;
assign i[11655]= 16'hf17;
assign i[11656]= 16'h1081;
assign i[11657]= 16'h1219;
assign i[11658]= 16'h13d9;
assign i[11659]= 16'h15ba;
assign i[11660]= 16'h17b4;
assign i[11661]= 16'h19bf;
assign i[11662]= 16'h1bd0;
assign i[11663]= 16'h1ddd;
assign i[11664]= 16'h1fda;
assign i[11665]= 16'h21bc;
assign i[11666]= 16'h2377;
assign i[11667]= 16'h2501;
assign i[11668]= 16'h264d;
assign i[11669]= 16'h2753;
assign i[11670]= 16'h2808;
assign i[11671]= 16'h2864;
assign i[11672]= 16'h2860;
assign i[11673]= 16'h27f7;
assign i[11674]= 16'h2724;
assign i[11675]= 16'h25e5;
assign i[11676]= 16'h2439;
assign i[11677]= 16'h221f;
assign i[11678]= 16'h1f9a;
assign i[11679]= 16'h1cae;
assign i[11680]= 16'h195f;
assign i[11681]= 16'h15b4;
assign i[11682]= 16'h11b6;
assign i[11683]= 16'hd6c;
assign i[11684]= 16'h8e3;
assign i[11685]= 16'h426;
assign i[11686]= 16'hff43;
assign i[11687]= 16'hfa46;
assign i[11688]= 16'hf542;
assign i[11689]= 16'hf045;
assign i[11690]= 16'heb61;
assign i[11691]= 16'he6a8;
assign i[11692]= 16'he22e;
assign i[11693]= 16'hde03;
assign i[11694]= 16'hda3c;
assign i[11695]= 16'hd6eb;
assign i[11696]= 16'hd420;
assign i[11697]= 16'hd1ed;
assign i[11698]= 16'hd060;
assign i[11699]= 16'hcf85;
assign i[11700]= 16'hcf65;
assign i[11701]= 16'hd009;
assign i[11702]= 16'hd173;
assign i[11703]= 16'hd3a2;
assign i[11704]= 16'hd692;
assign i[11705]= 16'hda39;
assign i[11706]= 16'hde8b;
assign i[11707]= 16'he375;
assign i[11708]= 16'he8e2;
assign i[11709]= 16'heeb7;
assign i[11710]= 16'hf4d8;
assign i[11711]= 16'hfb25;
assign i[11712]= 16'h17b;
assign i[11713]= 16'h7b9;
assign i[11714]= 16'hdba;
assign i[11715]= 16'h135d;
assign i[11716]= 16'h1880;
assign i[11717]= 16'h1d05;
assign i[11718]= 16'h20d3;
assign i[11719]= 16'h23d3;
assign i[11720]= 16'h25f5;
assign i[11721]= 16'h272e;
assign i[11722]= 16'h277a;
assign i[11723]= 16'h26db;
assign i[11724]= 16'h255a;
assign i[11725]= 16'h2307;
assign i[11726]= 16'h1ff5;
assign i[11727]= 16'h1c3e;
assign i[11728]= 16'h1802;
assign i[11729]= 16'h1361;
assign i[11730]= 16'he80;
assign i[11731]= 16'h982;
assign i[11732]= 16'h48d;
assign i[11733]= 16'hffc4;
assign i[11734]= 16'hfb44;
assign i[11735]= 16'hf72c;
assign i[11736]= 16'hf392;
assign i[11737]= 16'hf088;
assign i[11738]= 16'hee1a;
assign i[11739]= 16'hec4c;
assign i[11740]= 16'heb1d;
assign i[11741]= 16'hea86;
assign i[11742]= 16'hea79;
assign i[11743]= 16'heae4;
assign i[11744]= 16'hebb1;
assign i[11745]= 16'hecc5;
assign i[11746]= 16'hee06;
assign i[11747]= 16'hef58;
assign i[11748]= 16'hf0a0;
assign i[11749]= 16'hf1c5;
assign i[11750]= 16'hf2b1;
assign i[11751]= 16'hf353;
assign i[11752]= 16'hf39f;
assign i[11753]= 16'hf38e;
assign i[11754]= 16'hf321;
assign i[11755]= 16'hf25c;
assign i[11756]= 16'hf14b;
assign i[11757]= 16'hf001;
assign i[11758]= 16'hee93;
assign i[11759]= 16'hed1a;
assign i[11760]= 16'hebb4;
assign i[11761]= 16'hea7e;
assign i[11762]= 16'he996;
assign i[11763]= 16'he918;
assign i[11764]= 16'he91d;
assign i[11765]= 16'he9ba;
assign i[11766]= 16'heaff;
assign i[11767]= 16'hecf6;
assign i[11768]= 16'hef9f;
assign i[11769]= 16'hf2f7;
assign i[11770]= 16'hf6f1;
assign i[11771]= 16'hfb78;
assign i[11772]= 16'h71;
assign i[11773]= 16'h5bc;
assign i[11774]= 16'hb34;
assign i[11775]= 16'h10af;
assign i[11776]= 16'h1601;
assign i[11777]= 16'h1afd;
assign i[11778]= 16'h1f7a;
assign i[11779]= 16'h234e;
assign i[11780]= 16'h2656;
assign i[11781]= 16'h2874;
assign i[11782]= 16'h298f;
assign i[11783]= 16'h2999;
assign i[11784]= 16'h288b;
assign i[11785]= 16'h2667;
assign i[11786]= 16'h2339;
assign i[11787]= 16'h1f16;
assign i[11788]= 16'h1a19;
assign i[11789]= 16'h1466;
assign i[11790]= 16'he28;
assign i[11791]= 16'h78e;
assign i[11792]= 16'hc8;
assign i[11793]= 16'hfa0d;
assign i[11794]= 16'hf38e;
assign i[11795]= 16'hed7d;
assign i[11796]= 16'he808;
assign i[11797]= 16'he359;
assign i[11798]= 16'hdf93;
assign i[11799]= 16'hdcd2;
assign i[11800]= 16'hdb29;
assign i[11801]= 16'hdaa4;
assign i[11802]= 16'hdb46;
assign i[11803]= 16'hdd08;
assign i[11804]= 16'hdfdd;
assign i[11805]= 16'he3ae;
assign i[11806]= 16'he860;
assign i[11807]= 16'hedcf;
assign i[11808]= 16'hf3d7;
assign i[11809]= 16'hfa4c;
assign i[11810]= 16'h104;
assign i[11811]= 16'h7d5;
assign i[11812]= 16'he92;
assign i[11813]= 16'h1513;
assign i[11814]= 16'h1b33;
assign i[11815]= 16'h20d0;
assign i[11816]= 16'h25ce;
assign i[11817]= 16'h2a14;
assign i[11818]= 16'h2d91;
assign i[11819]= 16'h3037;
assign i[11820]= 16'h3200;
assign i[11821]= 16'h32eb;
assign i[11822]= 16'h32f8;
assign i[11823]= 16'h3231;
assign i[11824]= 16'h309f;
assign i[11825]= 16'h2e51;
assign i[11826]= 16'h2b57;
assign i[11827]= 16'h27c5;
assign i[11828]= 16'h23ad;
assign i[11829]= 16'h1f26;
assign i[11830]= 16'h1a42;
assign i[11831]= 16'h1519;
assign i[11832]= 16'hfbe;
assign i[11833]= 16'ha47;
assign i[11834]= 16'h4c7;
assign i[11835]= 16'hff53;
assign i[11836]= 16'hf9fa;
assign i[11837]= 16'hf4d0;
assign i[11838]= 16'hefe6;
assign i[11839]= 16'heb4c;
assign i[11840]= 16'he711;
assign i[11841]= 16'he344;
assign i[11842]= 16'hdff3;
assign i[11843]= 16'hdd29;
assign i[11844]= 16'hdaf0;
assign i[11845]= 16'hd951;
assign i[11846]= 16'hd852;
assign i[11847]= 16'hd7f8;
assign i[11848]= 16'hd843;
assign i[11849]= 16'hd931;
assign i[11850]= 16'hdabe;
assign i[11851]= 16'hdce0;
assign i[11852]= 16'hdf8b;
assign i[11853]= 16'he2b1;
assign i[11854]= 16'he63e;
assign i[11855]= 16'hea1f;
assign i[11856]= 16'hee3c;
assign i[11857]= 16'hf27b;
assign i[11858]= 16'hf6c3;
assign i[11859]= 16'hfafb;
assign i[11860]= 16'hff08;
assign i[11861]= 16'h2d4;
assign i[11862]= 16'h649;
assign i[11863]= 16'h957;
assign i[11864]= 16'hbee;
assign i[11865]= 16'he05;
assign i[11866]= 16'hf99;
assign i[11867]= 16'h10aa;
assign i[11868]= 16'h113e;
assign i[11869]= 16'h1161;
assign i[11870]= 16'h1122;
assign i[11871]= 16'h1096;
assign i[11872]= 16'hfd4;
assign i[11873]= 16'hef5;
assign i[11874]= 16'he15;
assign i[11875]= 16'hd4f;
assign i[11876]= 16'hcbc;
assign i[11877]= 16'hc74;
assign i[11878]= 16'hc8b;
assign i[11879]= 16'hd11;
assign i[11880]= 16'he0f;
assign i[11881]= 16'hf8a;
assign i[11882]= 16'h117f;
assign i[11883]= 16'h13e5;
assign i[11884]= 16'h16ad;
assign i[11885]= 16'h19c1;
assign i[11886]= 16'h1d06;
assign i[11887]= 16'h205c;
assign i[11888]= 16'h23a1;
assign i[11889]= 16'h26af;
assign i[11890]= 16'h2962;
assign i[11891]= 16'h2b95;
assign i[11892]= 16'h2d27;
assign i[11893]= 16'h2df9;
assign i[11894]= 16'h2df5;
assign i[11895]= 16'h2d07;
assign i[11896]= 16'h2b27;
assign i[11897]= 16'h2853;
assign i[11898]= 16'h2490;
assign i[11899]= 16'h1fef;
assign i[11900]= 16'h1a88;
assign i[11901]= 16'h1479;
assign i[11902]= 16'hdea;
assign i[11903]= 16'h704;
assign i[11904]= 16'hfff9;
assign i[11905]= 16'hf8f9;
assign i[11906]= 16'hf236;
assign i[11907]= 16'hebe2;
assign i[11908]= 16'he62b;
assign i[11909]= 16'he139;
assign i[11910]= 16'hdd2f;
assign i[11911]= 16'hda29;
assign i[11912]= 16'hd838;
assign i[11913]= 16'hd765;
assign i[11914]= 16'hd7b0;
assign i[11915]= 16'hd90e;
assign i[11916]= 16'hdb6b;
assign i[11917]= 16'hdeaa;
assign i[11918]= 16'he2a6;
assign i[11919]= 16'he736;
assign i[11920]= 16'hec29;
assign i[11921]= 16'hf14e;
assign i[11922]= 16'hf672;
assign i[11923]= 16'hfb60;
assign i[11924]= 16'hffea;
assign i[11925]= 16'h3e3;
assign i[11926]= 16'h728;
assign i[11927]= 16'h997;
assign i[11928]= 16'hb1d;
assign i[11929]= 16'hbaa;
assign i[11930]= 16'hb3b;
assign i[11931]= 16'h9d5;
assign i[11932]= 16'h787;
assign i[11933]= 16'h466;
assign i[11934]= 16'h91;
assign i[11935]= 16'hfc2c;
assign i[11936]= 16'hf75d;
assign i[11937]= 16'hf251;
assign i[11938]= 16'hed34;
assign i[11939]= 16'he832;
assign i[11940]= 16'he374;
assign i[11941]= 16'hdf21;
assign i[11942]= 16'hdb5a;
assign i[11943]= 16'hd839;
assign i[11944]= 16'hd5d3;
assign i[11945]= 16'hd434;
assign i[11946]= 16'hd361;
assign i[11947]= 16'hd356;
assign i[11948]= 16'hd408;
assign i[11949]= 16'hd566;
assign i[11950]= 16'hd757;
assign i[11951]= 16'hd9c1;
assign i[11952]= 16'hdc81;
assign i[11953]= 16'hdf77;
assign i[11954]= 16'he27f;
assign i[11955]= 16'he577;
assign i[11956]= 16'he83d;
assign i[11957]= 16'heab4;
assign i[11958]= 16'hecc4;
assign i[11959]= 16'hee57;
assign i[11960]= 16'hef60;
assign i[11961]= 16'hefd6;
assign i[11962]= 16'hefb6;
assign i[11963]= 16'hef06;
assign i[11964]= 16'hedce;
assign i[11965]= 16'hec1d;
assign i[11966]= 16'hea07;
assign i[11967]= 16'he7a4;
assign i[11968]= 16'he50b;
assign i[11969]= 16'he25a;
assign i[11970]= 16'hdfa9;
assign i[11971]= 16'hdd16;
assign i[11972]= 16'hdab7;
assign i[11973]= 16'hd8a3;
assign i[11974]= 16'hd6ee;
assign i[11975]= 16'hd5a6;
assign i[11976]= 16'hd4d4;
assign i[11977]= 16'hd480;
assign i[11978]= 16'hd4a9;
assign i[11979]= 16'hd54c;
assign i[11980]= 16'hd661;
assign i[11981]= 16'hd7dc;
assign i[11982]= 16'hd9af;
assign i[11983]= 16'hdbc6;
assign i[11984]= 16'hde0f;
assign i[11985]= 16'he075;
assign i[11986]= 16'he2e2;
assign i[11987]= 16'he543;
assign i[11988]= 16'he782;
assign i[11989]= 16'he98f;
assign i[11990]= 16'heb59;
assign i[11991]= 16'hecd3;
assign i[11992]= 16'hedf2;
assign i[11993]= 16'heeae;
assign i[11994]= 16'hef04;
assign i[11995]= 16'heef2;
assign i[11996]= 16'hee79;
assign i[11997]= 16'hed9c;
assign i[11998]= 16'hec63;
assign i[11999]= 16'head4;
assign i[12000]= 16'he8fa;
assign i[12001]= 16'he6e0;
assign i[12002]= 16'he492;
assign i[12003]= 16'he21b;
assign i[12004]= 16'hdf8a;
assign i[12005]= 16'hdcea;
assign i[12006]= 16'hda48;
assign i[12007]= 16'hd7b1;
assign i[12008]= 16'hd530;
assign i[12009]= 16'hd2d0;
assign i[12010]= 16'hd09c;
assign i[12011]= 16'hce9f;
assign i[12012]= 16'hcce1;
assign i[12013]= 16'hcb6b;
assign i[12014]= 16'hca45;
assign i[12015]= 16'hc977;
assign i[12016]= 16'hc906;
assign i[12017]= 16'hc8f8;
assign i[12018]= 16'hc952;
assign i[12019]= 16'hca16;
assign i[12020]= 16'hcb46;
assign i[12021]= 16'hcce2;
assign i[12022]= 16'hcee9;
assign i[12023]= 16'hd157;
assign i[12024]= 16'hd427;
assign i[12025]= 16'hd752;
assign i[12026]= 16'hdacd;
assign i[12027]= 16'hde8d;
assign i[12028]= 16'he284;
assign i[12029]= 16'he6a4;
assign i[12030]= 16'heada;
assign i[12031]= 16'hef16;
assign i[12032]= 16'hf343;
assign i[12033]= 16'hf74f;
assign i[12034]= 16'hfb26;
assign i[12035]= 16'hfeb6;
assign i[12036]= 16'h1ed;
assign i[12037]= 16'h4bd;
assign i[12038]= 16'h719;
assign i[12039]= 16'h8f6;
assign i[12040]= 16'ha4e;
assign i[12041]= 16'hb1c;
assign i[12042]= 16'hb61;
assign i[12043]= 16'hb21;
assign i[12044]= 16'ha63;
assign i[12045]= 16'h934;
assign i[12046]= 16'h7a1;
assign i[12047]= 16'h5bb;
assign i[12048]= 16'h396;
assign i[12049]= 16'h149;
assign i[12050]= 16'hfee9;
assign i[12051]= 16'hfc8b;
assign i[12052]= 16'hfa47;
assign i[12053]= 16'hf832;
assign i[12054]= 16'hf65f;
assign i[12055]= 16'hf4df;
assign i[12056]= 16'hf3bf;
assign i[12057]= 16'hf30b;
assign i[12058]= 16'hf2c7;
assign i[12059]= 16'hf2f9;
assign i[12060]= 16'hf39d;
assign i[12061]= 16'hf4b0;
assign i[12062]= 16'hf62a;
assign i[12063]= 16'hf7fe;
assign i[12064]= 16'hfa1e;
assign i[12065]= 16'hfc7b;
assign i[12066]= 16'hff02;
assign i[12067]= 16'h1a0;
assign i[12068]= 16'h445;
assign i[12069]= 16'h6de;
assign i[12070]= 16'h959;
assign i[12071]= 16'hba7;
assign i[12072]= 16'hdbd;
assign i[12073]= 16'hf8f;
assign i[12074]= 16'h1115;
assign i[12075]= 16'h124c;
assign i[12076]= 16'h1332;
assign i[12077]= 16'h13c7;
assign i[12078]= 16'h1410;
assign i[12079]= 16'h1413;
assign i[12080]= 16'h13d8;
assign i[12081]= 16'h1369;
assign i[12082]= 16'h12d0;
assign i[12083]= 16'h1218;
assign i[12084]= 16'h114c;
assign i[12085]= 16'h1078;
assign i[12086]= 16'hfa5;
assign i[12087]= 16'hedc;
assign i[12088]= 16'he26;
assign i[12089]= 16'hd87;
assign i[12090]= 16'hd04;
assign i[12091]= 16'hca0;
assign i[12092]= 16'hc5d;
assign i[12093]= 16'hc3b;
assign i[12094]= 16'hc38;
assign i[12095]= 16'hc53;
assign i[12096]= 16'hc89;
assign i[12097]= 16'hcd7;
assign i[12098]= 16'hd3b;
assign i[12099]= 16'hdb2;
assign i[12100]= 16'he3b;
assign i[12101]= 16'hed4;
assign i[12102]= 16'hf7d;
assign i[12103]= 16'h1036;
assign i[12104]= 16'h1101;
assign i[12105]= 16'h11de;
assign i[12106]= 16'h12d1;
assign i[12107]= 16'h13dd;
assign i[12108]= 16'h1503;
assign i[12109]= 16'h1647;
assign i[12110]= 16'h17ab;
assign i[12111]= 16'h1930;
assign i[12112]= 16'h1ad6;
assign i[12113]= 16'h1c9d;
assign i[12114]= 16'h1e82;
assign i[12115]= 16'h2083;
assign i[12116]= 16'h2299;
assign i[12117]= 16'h24bf;
assign i[12118]= 16'h26ed;
assign i[12119]= 16'h2919;
assign i[12120]= 16'h2b3a;
assign i[12121]= 16'h2d45;
assign i[12122]= 16'h2f2e;
assign i[12123]= 16'h30ec;
assign i[12124]= 16'h3272;
assign i[12125]= 16'h33b5;
assign i[12126]= 16'h34ad;
assign i[12127]= 16'h3551;
assign i[12128]= 16'h3598;
assign i[12129]= 16'h357d;
assign i[12130]= 16'h34fc;
assign i[12131]= 16'h3410;
assign i[12132]= 16'h32b9;
assign i[12133]= 16'h30f5;
assign i[12134]= 16'h2ec8;
assign i[12135]= 16'h2c32;
assign i[12136]= 16'h2938;
assign i[12137]= 16'h25de;
assign i[12138]= 16'h222a;
assign i[12139]= 16'h1e22;
assign i[12140]= 16'h19cd;
assign i[12141]= 16'h1531;
assign i[12142]= 16'h1058;
assign i[12143]= 16'hb48;
assign i[12144]= 16'h60b;
assign i[12145]= 16'haa;
assign i[12146]= 16'hfb31;
assign i[12147]= 16'hf5a7;
assign i[12148]= 16'hf01a;
assign i[12149]= 16'hea96;
assign i[12150]= 16'he529;
assign i[12151]= 16'hdfe1;
assign i[12152]= 16'hdacd;
assign i[12153]= 16'hd5fd;
assign i[12154]= 16'hd183;
assign i[12155]= 16'hcd70;
assign i[12156]= 16'hc9d4;
assign i[12157]= 16'hc6c0;
assign i[12158]= 16'hc445;
assign i[12159]= 16'hc272;
assign i[12160]= 16'hc152;
assign i[12161]= 16'hc0f3;
assign i[12162]= 16'hc15a;
assign i[12163]= 16'hc28e;
assign i[12164]= 16'hc48f;
assign i[12165]= 16'hc75a;
assign i[12166]= 16'hcae9;
assign i[12167]= 16'hcf2f;
assign i[12168]= 16'hd41e;
assign i[12169]= 16'hd9a2;
assign i[12170]= 16'hdfa2;
assign i[12171]= 16'he605;
assign i[12172]= 16'hecaa;
assign i[12173]= 16'hf374;
assign i[12174]= 16'hfa3e;
assign i[12175]= 16'he7;
assign i[12176]= 16'h74c;
assign i[12177]= 16'hd4d;
assign i[12178]= 16'h12ca;
assign i[12179]= 16'h17a5;
assign i[12180]= 16'h1bc5;
assign i[12181]= 16'h1f16;
assign i[12182]= 16'h2185;
assign i[12183]= 16'h2309;
assign i[12184]= 16'h239a;
assign i[12185]= 16'h2337;
assign i[12186]= 16'h21e6;
assign i[12187]= 16'h1fb0;
assign i[12188]= 16'h1ca3;
assign i[12189]= 16'h18d3;
assign i[12190]= 16'h1457;
assign i[12191]= 16'hf49;
assign i[12192]= 16'h9c6;
assign i[12193]= 16'h3ed;
assign i[12194]= 16'hfddf;
assign i[12195]= 16'hf7ba;
assign i[12196]= 16'hf19e;
assign i[12197]= 16'hebac;
assign i[12198]= 16'he600;
assign i[12199]= 16'he0b6;
assign i[12200]= 16'hdbe7;
assign i[12201]= 16'hd7a9;
assign i[12202]= 16'hd40e;
assign i[12203]= 16'hd127;
assign i[12204]= 16'hcf00;
assign i[12205]= 16'hcda1;
assign i[12206]= 16'hcd10;
assign i[12207]= 16'hcd4e;
assign i[12208]= 16'hce5a;
assign i[12209]= 16'hd02f;
assign i[12210]= 16'hd2c5;
assign i[12211]= 16'hd611;
assign i[12212]= 16'hda05;
assign i[12213]= 16'hde90;
assign i[12214]= 16'he3a0;
assign i[12215]= 16'he91f;
assign i[12216]= 16'heef5;
assign i[12217]= 16'hf509;
assign i[12218]= 16'hfb41;
assign i[12219]= 16'h17f;
assign i[12220]= 16'h7a9;
assign i[12221]= 16'hda1;
assign i[12222]= 16'h1349;
assign i[12223]= 16'h1886;
assign i[12224]= 16'h1d3c;
assign i[12225]= 16'h2153;
assign i[12226]= 16'h24b4;
assign i[12227]= 16'h274d;
assign i[12228]= 16'h290c;
assign i[12229]= 16'h29e8;
assign i[12230]= 16'h29da;
assign i[12231]= 16'h28df;
assign i[12232]= 16'h26fd;
assign i[12233]= 16'h243b;
assign i[12234]= 16'h20aa;
assign i[12235]= 16'h1c5d;
assign i[12236]= 16'h176c;
assign i[12237]= 16'h11f6;
assign i[12238]= 16'hc1a;
assign i[12239]= 16'h5fd;
assign i[12240]= 16'hffc5;
assign i[12241]= 16'hf997;
assign i[12242]= 16'hf39b;
assign i[12243]= 16'hedf5;
assign i[12244]= 16'he8c9;
assign i[12245]= 16'he437;
assign i[12246]= 16'he05a;
assign i[12247]= 16'hdd47;
assign i[12248]= 16'hdb11;
assign i[12249]= 16'hd9c0;
assign i[12250]= 16'hd959;
assign i[12251]= 16'hd9d8;
assign i[12252]= 16'hdb35;
assign i[12253]= 16'hdd5f;
assign i[12254]= 16'he042;
assign i[12255]= 16'he3c3;
assign i[12256]= 16'he7c4;
assign i[12257]= 16'hec24;
assign i[12258]= 16'hf0bf;
assign i[12259]= 16'hf573;
assign i[12260]= 16'hfa1a;
assign i[12261]= 16'hfe94;
assign i[12262]= 16'h2bf;
assign i[12263]= 16'h680;
assign i[12264]= 16'h9bf;
assign i[12265]= 16'hc67;
assign i[12266]= 16'he6b;
assign i[12267]= 16'hfbf;
assign i[12268]= 16'h1062;
assign i[12269]= 16'h1053;
assign i[12270]= 16'hf99;
assign i[12271]= 16'he3f;
assign i[12272]= 16'hc53;
assign i[12273]= 16'h9e6;
assign i[12274]= 16'h70d;
assign i[12275]= 16'h3dd;
assign i[12276]= 16'h6b;
assign i[12277]= 16'hfccf;
assign i[12278]= 16'hf91c;
assign i[12279]= 16'hf567;
assign i[12280]= 16'hf1c2;
assign i[12281]= 16'hee3d;
assign i[12282]= 16'heae4;
assign i[12283]= 16'he7c3;
assign i[12284]= 16'he4e1;
assign i[12285]= 16'he243;
assign i[12286]= 16'hdfeb;
assign i[12287]= 16'hddda;
